��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��33�z_�`�f����EW^7"q5���K��Ҋ���CU��ˑ�v~,�ynfP\��j��I�qS�of�*͐v�C��ڋ�I�3�f���e"���m�Dm��	�ӍE��O����/
�=2�rU�&��07���eև�`�vr�M�q�.,+�`����-\���'�]��ڙ�WT�5��3���d��� ���WTlc��E���v��̌�A$���	�+n+Y��rU�@X��rH�Ze"\pq2^Ԁ\�/4�d�O�X7��2����XجH�/�y$�1@agCGY�Yg\�(<%��I�6��6��^�6;�;s��������[qqX�$�+TևeC���T��ّ��P�iwk��n�0�Z�!f���S�4�5����G��2�/�dj_z�j�SC�(��I�`����l�����c��G��gk�����dBm�n�*e�[�9똢h9�.�t�ꋝ��@ۭ֝O�}�1>w�t�'���qS�7�C�r���_�M=����IB�c��#�����|ҸG^��2�g�D���)�|~s�o;��q�k6L'T��&�����
A�������i��V_��!�V~�yW�<��T��vB��:�>r
�xv vd0AL h&B�}X���L�dH
(���(����������M�:�q%�����;�~|�"M�]��#�X��p/���B�E��~�$���b{��(�OM*6�s��e~QelHC��(��y��=�]W<�ۘ���[�	>-�� |���r��Mn�Y���eP��]���R"��!~�u"?$Z1�� D��g$�ԚFӞ6I,��zT܍ݙ7V,9�$�J��	��k_��%�PQ��I����|G���Es�"����>"�gΏ���7|Y�zXF�V�P��+��R.-c��:X���󟵱N��1�S|'��mU)���p�d8�{2�\Ů��5zC��4�R(B����Ə�8��X��Q;�f�K��6�3��c�ӥ�<���2.�|F���#Nr�����˕�ND�����}�UJ�iD����R 1�' �9o�*��Tj��h����Z@l�l�x9�͗I=>�EM/�:�)�]���6�;>o}���*�5� �$_�EK��+}dl��%)U.����֨�u��U����o�lm ][Rg��44��^^�+��O�`H[�i�M����4-L�)��S��bY�Z�Lt:�v�F���N��46�z�l�d��+P%��ӭb�ǋ�y'K�Y�6`�GI!
>0�OI�B��Z&��;���3����!�*�C���͍G�b��;E|���8�VO-�Ռ��$�?N��OeHW��;iS�����H�َ���U'�I�z|s�2�24��
Ɨ�o[]@�Z���S5oz�g��1R)�c0�����1w
ܫ��V3	�N�r�s\�ǥ�$L��f�¸�]�H�6���NհO�4��O������3yo��zCd�Wi�\C�&��8w{�'�̢yn�pH.7:�¼�o�a��ۥ�b�V!�eQ-�l�{�Ι"���)W���?�tr�#���������y�u⟬�3���%be��	���|γ�L�����A���hP�w�#��>�e%-$���1����EQg�E����!/�0LA�<��-F�u��f��s-�a0=[h�D���o�l~Mh�N��Έ�8�4�t,��=p�[�:�S#�?O L�;�sY4�G�RI�o)r:�Q,B�����w�R6dkr��NW;!8���Iue���Dn�i���QZ���e?;�츆����<��:K.g���݁��n���p1جE'3�5-�L|�O6P#ָ֚�v�}�b~8T_�@-�捯�Rr���-,��,�c���o,`���v��O�5xHe���n�A��!W�~7��|��C�������n��"� Z�wB�T�1&_�י���UeQ���_O��|X���9�q	��,)Z��!���,�r�OB�Y;�Z$1U���秷����+�i�"���H8_}�Q��k������e8������L��E?�������`�c�u�ד� ��]w��◯2��P;7��i�}��v��PO�ӭ�T�p	�!ygia�%ȎY����Qc�ƥ�)��?���������R�ɬӊ��j]ő޹,n�+|)F�.q�GM�v����lȝ�l�Q��wR����sY"vv���������]Y;l�d)u��2���/aOÃ��/��6e�A�K)�>]�2K	�3�&@W�?]͌�`�:�&���C�Rۘ�ew��'~U�^����ee
��e�I��.˥/AM�4��{!�DbT�
`6��Tgސps<B$&(�7��t�%Y�/���sz�/B���p����9��� Ʀ~gm�汌����$�nS��V���8C}�wd���\���	��-��
Mb���`	wlw
�*?wiT�r��c5C�a�J�f�ǨO��f
.�áwK����7W�X��E�.�;ʼ�YO~˔�����{ݲb=��8-�x�k�4�>�9�ũiTw��E�2��j�XYT���q�!*L1�2����(�YJ>$?.Q�y)m��]���<��K8�)g�t"Ƒly=g
j(�.�}�?qC��k�
W�)��V�:��[�&��3���N�����cg�,���Cd¯0s��^�G��:
�Wәk:�$>�����>%n�aoM~�.�3�)��Ԛ��43
^/� ���l��u8�~��#��b�0e�́/&N7�	�ζg��U��_#�y& '`��qƴ�;c�,D*���Oo���ٕ�����O���{���	�_=&P��D�Լ��ޒB܇M4I�D��|;g$ɥ�̅ms(��ָ�1xNl�h�2�K\�W�SU:B~��2���E(q�jrxr�*4"�߲glڻ9j�-Ǳ�Z�w r�p?6��eN���7K�K4
.;�kMm�M����s��Qey�2����y��F���ռL�-FM�"��>fC��塍5/����������	��a�:���((:��u6��qT�+Jґ?i�S�-d�Ór*����{ݒ�[���A�ؒ�o�����f(m��3�h�$�l>m�0��Y����A-�4�3����]���,~�Ƹ���ɑ����=�F6է�mo���`� �-wj
����������锌�v���J�3��(b/Cj}9��R��O�4qk�P=�rm���(zɬ��S˓�-�Ĩ�d�&��ז����	���Ea�F�ME���IVaBZ6=нSJ0��za�.�<J�	�h�_i�������Hۻ�ۏrF%�=FD����,tv���޻��
��4.Wn�J����:��a����6�%\�k�	9�n�0 �n%V��@yu{L���޸��x����l�	�����P����O"n�Ų�;�A�h�qlT��\n-��K��Njz��#��UA>���S�KT�Rā��Ga�FIڳ�]B��\T�fZ���D���c�m�Y�BlSQh0���(Gz8ew�HuwT��o�R�����2Q#���y	�$�78�G�<gu�K�S�k^
QX�DrsGff�8D���A�ײ]5��Ƚ��55��^��;h���o\���Kz���	,4Ŋ�E�?\�Aι�2yv#�U7b�����|3L�~���K$A�7R+�KQ;�~�]�f������R�h"l��9����
6=����P������v��4�	������J�Mk<��8���G(Iu���f������-��x�H?��pʭQ�lV���h�#|�G��˛���8��fͰ���<���	rU�h-_�W�(ӏ�(�X��w��+<[�ΐe{�qE��'B��Eiv�ȍF�:@���ϰ���6��"+J�n��òwc[]��
&%���e��R�d�K'���x�5AݜnVԜ����5���&ڡb�D}M�0���-�D	���خ��o�F@�t��I�g'�+oQ�c�L�Ȭ���e�,L�E�y�t�y�
�+Ւ�ۓ@ˋ�dL�⹔r�L�8�r	X�� l��^�J����Ȝ����g+>T��#^�]���,ۈ�[O��yԥ.=I��ҭ đzK��Ar��J�C�7m�j�TY�H�r\��N��n�jj��~�Q��3�otovi%1��Q	�o��̸M���X�n�'�?o����3h%�J��P�a7a�A!�\-%���;�@������u7������`�(�u��)t*}�C9��6�(S���w��0)�:�^��aW���S�^��!␚���;U���`я��b9���r�{�S��[պU�:�2η)���%}��6��K4��
$�tu�cx����8I?��?7 ���n{'*��SWW�%�����E�t֠����N�a�y��'��蔓BB�<h�Vd0R�\�~!�܊\��(�yT�A��C�ֺl9u�;O�Wށfp�C�)�l4��]��yD�&M�]D�`M�!_t�N� �m��m���0�dHA�r#u����l�Ga��Cъ����f!+�+�XE�ayvj$*�jbۛ=���q�����	X~�m�͌�6�����	�����xg9d؅n=Ŧx��!h��mT���7��$�AdZ�	Q^gS�o+�Q�sS�~��t��D<y��ә�
5ZX׷:b	�?�#�����OW�5�I$��8�o��L��E�&-�d ���$F8M5[ G/�^��ģ�rb��F��Ӟz�^�C<h���?��/���	�� �,٧�Tێ� 6A?�J��"x�.:���$�d��D[ΙK��W�lq*\�R��pvq�(��0���]4ԓ���'��Mc$��WI�(��k#�+��S+t?}���\��{��?}�����U��>�PcɆ3jYMhF}��Qcbԉ������Hb�������p}L�L�Z�ޓ�鈒 �AusM}p��[���
G,�tƪC�%�9<{-��l�7�O�DrQ��x�O���Oyq��7;e��9�5Z��?a��1��|��w��*t#��! 	�-[�h nS~ATe���H�Y�N�Y�\��ְ�011n�4�����m��W���h�nB6B������*���^�!'�k�%�jQ�e��v�\�\�Veo�q���C��fh؀�����V`B�5ڄ.�(���߈i��C7�$�MO��8�{��Ƶ̴������G��.2��Y}�y��T�րq]��F��"�V,E4̖m�OR���~���8A�d���^h9���,:�X��O���i��~y�c�I�P�[[r��)	�1��w�������
����O��/d3:���u1u�27���]��Y����3ހC0�c�{�g�~�=��Ľ揪�Tx�;���W&���x/<[��.�����y\���'aR�
�
"��s�s��nm�R��ۄ�A��������>g�śn��f0ځ��LnUY�yw��zoա.Y��U��|}��T~��L��D&]I��1yt�ߊ>K��{A5����CWEi����� ���ΐۼ�=�A"d�fc���p��>�����q�K�Ř�9$l�M
[/�2�=���Ao�jo�mg��;�\�Ɍ��}�i<I����҆�S���4��$�;A�/!u�V}}<k�X_�I�������)�7�،�X�S�߬{%]�R��b�����������S	.�3���?|���"�	|mb���t���ɕ�5_W=��eμ��|*Dz�fU�S+%���O�3M_��t	����4"�:�����W���(�N����@�-(]�Φ����2{�����/%V�RBf��p"��إ�ؕL�£Mnqt���n�̶�	,�8w�`�d8���J��4&�g�JpP�?b�-�/Sf���bC|5�3���xaJ�2�� ���t� 6ٔ1�S|Ynsw�;?6���Kw�I�Zq�{��H�!O��*4��9b�V�P��B��b�����Q�"�и�ĸ����Ce�B��<-��Z���3^�F,
��4R����iՌ��`9��a3d�Tbx���%�ǀ��[�v�9SهӬ����nN�s�er��w��C=V���Z7:7��O1C�pp����s��t!#b���� �S�=��R��M��]+���F������𬆔���D��Ӱ�9������zS)��M�w��fPf����C�U>l2s3�?�9k%�Y�_��������I"cV��`�-'�Oſ�bz����u9=�2�r��9'�����{�#S����h�fWj�	{������CB��}\A}��l�y]%@�#J�f?��Yt��x�Q|.��&��j����=��1���-��G}���`=��!�+K�p�?ʄ�A�G��gm-��B	s�q6ٲ�����8���ͩ��]XT7����8��E�m9��@)�m�e2)�JF��U����rږ�b|�<���!e�ME�M��M�e���I�p@��r��Kjch��U�|{����vd�d��ծj������Rz-�8��m8u�MW-&<�F�A�?���^�+����QpA�Q�ק�2"�>5U���`�=iN�PX6 �ؔ�N�H}�ŗ|H��zNX�!�ݕ>E .�ss����9�z�Ȉ����^Þ���s3o��d�'Q���#��w��"�������*�W#���L|�����p|H�ؽi�x0��܍�sK�� ����)��� �p5�����R���ֹ�4�9�~���]�U�Jbo��\
7�	��h��7FG��OftEۃ��3�u�=b�]U��G�j!��t�������%J d�BVI���D��tB��d̴��蜔��+�b����Q�ߥ�Uٍ���f��W�(�z&4ۺu�K]�eqG��`���uĆ�^6''����]H�Xc�nj��,�١��'w@#�~U�+��ѹ����Z�+��8r��&�.��η��%�5O�cU���;*��Fh��d~Թ�m�v�� {�l	r�V��ʜQ�~�2\��fY��8�od�-D�{�u�ף����0T-^��	8#�Gl]j"6�۷0�K�yx�h�)�c97'�5.f�,��d���j����սJ�+�6k��*�^���Ku^[ib��EVG)�>��˓˛2n�^�\-{��n�;�a�n�����?Q�a:N7��lkh��f��,|YC�y/�EӉ[&>Fݝj�/�eh���0�=N�����"��-��;��B3SC]G�Yk�&��@�)VDW��m;a�5�}���
jAa�<%�	o�:����I�h�>�v�"�W�����g��&�v	x4)��}��l��nG�H4������c��j����L���2.:X̼�gfF3�[Mv%�:����<����g����D-�Ŋý�	V;�4���%��7���!�~V��B�c`����C�o�hmH<��_�� c� �ة0Ju�Z`�W�߫G[��(t�I���f��rȩ�X��C��+%lVϿ��#S�(���)h`�f��SI5�$	�W>�J�KZB�h�fu\ͱ#���qh�/Q
��=�/\d� (R����^1l�s�1��Oc���W���'���ENӴ�F�I9RjX�W)��Vz*lC�P��Xo�g�օ����'�^x��Zq�^'3�r�M�Q�P8g�p��4G�Ȅ�G1@`]	���Rz� ���;��Րs�i �8ɽ�R}�sY���h���}�1h[mj~ ��A�̭ĪQG� VN����Kbn�T��ԥ|���*�zՁMf��@�6��vv��[0@$)/]�#Ӧ:��z�7�Zm A.�(�(�U����+@J�z?ܢ,���☄7�#Aq�-kJZ�fH>zV+y�x�x*�?�"{b��W����V#���~��4W��BFH<*�v�\!�������̮�j�Zxj��D�_�~�(���ϐ��F1��C�����##�|ʪ���.�a(Z{we9낰Q��8.#tM���% u��f�S�99��FQX�T��:.&�N�?�. �k3pa&N�g1�	�������&B�a]W��6+qM��\��:��
���������{�(XZbO$ɠ\a0�@��j�[.�fw��R����(11�\W�J�7��U���w���_l;��&��J�٠2�:p0�;%Ln%�(t{">F��J����s�k�6�S7/�/��f�"�t8�x�UkCA��QᵀV��u_:��G�ֺ�Њ�zc�z79��m#�7�]<������E8���oE��㍡%�-�U���f���i�,!���a�+s� Q��j�#�m��`+�ar�*�uĔρ��4�`+$l)2x&�����2$<6���HBRp�+��r&��b�$%Q���5;-x�;!֢�,�\$���I�j�q�Q���g.���W�aJj,O�z�����H.�An��d�/iWo-����*�|�+E��W�<���zcg[�QZdr#�&�ղ){��՛�7����Ѭ,jh�nV��X��u8�s�A��k�oNXV��������:3y�G�r��c���Ç�%��\�;zLc�.�1 �"��3�����y�pj����
k��ֿ�$vAd2R�u��|�-h�ңD#�<���#Ɔ�`��2�!�����g���M�����D�X��H���_roL�&z1=L1ij*$�# _ε��L[���Ae-������t�/�D��-�$锥S�����/��g V�C�{�Pw��[�Q���0&�Ce��Qum4[h��{��6�ssI�T1^��M��e��T���1��N�M���ֽt��1J|i���W%H�Y4f?W�q�@���u�<��7'5]OZ�xO��&��Ŧ_��#:x�O��{��a��S~�uȏ�u}}��2�mwg'p�j�o4A�ow��N_��g�؈�a/�gE�Hߒn<�џ��!w[i���T&��u��q�3�w��q��=��mގ>�~�����)�I˔H"5��p�(k�]��l�8�֏qs�q
DK�3q�E(�x_��FA��0��B(k�Y{a?�&o��~�\S���GX(�-
�@�Nnil�؛+��0^Rm���E��G����^6���[�$�򉋛K;P�4�������ݰ��ӺV�Re�A�&�RC/!p<F#Bx�#;_�&����xn:e��7V���9�;KR�qC�oqt:wx��x�u2L�~��XsKf�!̠�hG	�:C>�XƟ�+U���}<��sFzLX�~'q�����9蛷]�aȥ��7�aT�8p�w�Q� �L>�;Zm���ĳ2m�&��H$s/��O�44J#����$�~�B�(]�h����D��9�B ����vm�\FzU1���Q9=��b�6�d�{n�nǱm	N��5��#:�V/�����W�6��| �%�>�TPM�c��E�z�1�~Lе�������Xy=��� �Cb��J�
j�S�
�#|9դ�YD!Nmy$�껶b*�"M&A����TxIv�}���v������u����BS��2���_��J�fn,���.�>�%��ᕵ~�{�y'��ğw�V=F�)
�w�J|3�7��c}����4R��|���d����Ȳ����fW�y����b�2��h!Y7�1{b츈I��[9�kA���Gm�e�ik�G�>��,���ǚ�c���(�S�^��`��{��@�
�eB	�a�%H��T��L%��b��a��FV�14c`�,�j�0��ά���i/���E\���Jqab����V���/4߳޷���ӺVėk��SLә֩���)ݓ��y�M��z�2�}���۝#��8?�C.n7�� �w_f �S�^|�6U���*���")���5�!�����8'��SÜb
��1���k ����lz=]�P�} 2Jt�S�d&�XOT���:ZW�TK���&:^n�u�5�
��:v�7O���}�����-�";v��|>��N2�f��x�6���D�`�<T��`/;�'�=^�
�Ģ��	|�:}��3}:�p�v􋊀	/��tw�+V
�GLO,���B߭�md��]T$3� �m������ ḓ���&�z�0;�u	J�r@{&#�D5�4��/;(#�h��ܟT�SK�2Y}�chE@�%�A�2��C�m �~ )�2#�� ��z�b�/Z�Y2�o��ݦc�pg`�CQE(4�+\T����eǬ�>�眸�O�=�
u*
_�3S��80�������;i����5Qs+�@�}j���[,��?���[6jbg�-���G�>_��I�����3���t�*U��,���Lr���9`�ݤo\�\��W�x��N�*��o�����ҭ�4  l��ibC��xf��otP��g���@�A�וG�j��{5+��3��S<+���G� �>!����=�q�Y$-����<��'KƻM\���XR �0�s�+;�z�!Ho.D�l��-�[.����ɵ�p [���@��Q�X�Y��>�xb8L�H����~����R�uD���ZqSO�u���� �\,f�c4�#��^�	ѫ��8z��:蒿��\�����"	М`>	�6%VU(2�!�Nq��0M�/S�L͢l��%g���}NL�Nc(�����sRZ�R����+��x���J��Yf��C�k�6c�7_X�Ȏ>"v��͕�٪�r��n~��ۣ�QP@ej�4�����_��z��$R��T�ʊ�{i�&��2����uY?+7w{S�6|���$f���/!��f��7��.�=��P�����Pr��;k��7�b�]����U��C8#~�n���%����q��I����4��Ш/�!؏�t�ڙ^ɓW79�q��@P85N���\���W�Œ2��킩�\�_��|V���\����T�	')�-}hB���%"�y�f��q*�a�'���V3v>6���Q˗b�J���V`��]D����N����}T�ku�����m��J�Q2ψ'���I��`"c����h�7ɑ,qd^�^@��K�Q�>M�k ֥vB�"��� F��0��+#�1���T6Tt8欲���U�xEz���D	z�e'�[�g
g���pM̗z���Ѷx�\��V¼�AOg4�&�ī��8)��Ⱥ|&�-TQyѮ���<�B�O��Y_l�I���8�W����=���u�9=���XL��mD.�2Ͷ̅?#ene����Yу)��O��A�(c��c��T��P��n��n_��j1,Ɩo���ڡ�K�Hn٧G���gXn%;"z,���LO����tSv��t�\	X�/j�Y��p�7Ʉ@oR��`<�p�Tq������J�~�7%]�,7��|Թ�7�f��0�9��i^<6�3�-�|c��*Ne]ku�����(e3<���+�,>{���	|���ي:k�T8]���~�9����<���ӳ©o|˃>�0Ѕ��Ie���2�l��XfB�C�u��y�O�4]j�N�oL��Kӻ	<�dU*��F����q�:���n����UO<RC�d�5!�r���F��6yR��yeu�Cӹ����|�����,�Q/q�QxU��|���7�Q��̼��K\��l-�0���.���}>�g�Q���=�͞���?�qy�M�w���d�I�p�W�u�>�ǧ���]�MA-,�bR�����26Ή�)q�MV'G��_���m���퇔�F_ �^0i`�~�Ć[��~�5�\{�r����<�e�Gk�3%Q̾�I���̳�p���*�B�+G�7)ޟ\�R����0����'�|#M��n�ZB~v���;Q<��%kJJpzE;&�
o���D{�vҠ���@ڳ��1_����-��
y��@p��bb�n�,��/MH~I	%�Y ���!����
�'g	���!���Hɰ'{
��[ȫ=�����I�Q��dW�}��uQ#��J��bv�!�N�Ϣr�=��4/��j�.r��K���㘪wDu�K�m�����˸�2.v�fI�t�Ǣ	K``��D�JOZ�
vA�E]���ԅ��.��Jy6Z�aӂ�Z�a��19�{Wu��v���>F�$�2R�)�Xd.C�<�#'�LJp����Z�Ҽۆ�wfVx�)|Z�ץ���`����⏜�H�}mƕ�{�Dס�x��� ċf]_�@c�v�*�o��{W��@#H�4��M��+����RX�y
ȋ���ͦ�n������o^��+��c8�)s3��y�z��]C�����X�)�9��6����^����M�����[����b��aG��(z��v G���8:9�
�����L�>� $B�U<cSJ�}���;������CK����7��GD�Ë&�-Ԧ�?�'�!�Ї	ߓ��A��z�hb�V�Q��dz�����M�a�?),���|��-��r�}iΝ�I-��!=�e�T�.b�����<3$h�9���R��:�+�Sos�����
l8��'�]F��k ��S��\~C�G�N�gr/������ׅ������<��{����@����1��	�!^FD�6�|�H(B"G4���Zg_RB�s��~ͻ��X����4m;Ȥ����Z���!��\6��X���I�3�Ͻ��,*�XQ
�f��mc�k���93l�N�S?ν1�A����!�r�nT��v���g!/�K��Dc2g�͆/�9����e�>y?��ȋ���M���O�|C�i.�h+��b�
�m2��98qw2���j��F�^�׶��ș���Zi�����)�y�H��X�*[pn)͟;}�:[1������:ޫw���^�x�>�[�d�Q��64��3}���̠���;؛�~�kk6�!�|�9ԟp/���c}�'�<�`G����a�E�!�f��DC����*B��M@%b���!���P����Ba�vq���U2���
`��-��=���Mb�U�`K�`���g�Һ��2��t�����a�ǸMu�������j?���|,�i�E<�rOkI~YG�X�q ,�K t�}�>Q�C�cv�9�v����n��%��OԶ9c�8�4a'!��Coq1L;�zy
��F1A$XԪ_����<���d *�vx͚�/�����"�_�:i��2�]P��0�/��7|4���ׯY6����b�4������?܍�gg%|=��思`�5�3OVU��F�|T��Nw|"h��DK1�l_b��ҽ�x[4c��Wk�_�hAd�0�<`�ΪA��w�{���%�R�]�O~m�c,k�%�E��7q�T�ͻ�XVI�����qe�A�"h�o�"��c-��3��n��r�AXAx���z��7Zj�I�������F��#�	R�g�kc��G�v�-��b�[�8�&�IK�Z0�$@���btz�@��H<���{�h�(��m�0�|��%��|��leb�G�p�eu���
�?���Է�:�d+�����1�G��lD������?�c�a�d�����4�Np#�:�P�č!+�*\&�يٓ���?�.�}Ȉ~/kվ�DY�ؤ _�9���#�y�4hf�����H��Ϣg�Q�����&!���q�/�o�X?5�b�FO�UCD�iPu�va��2��ڊ�oZ�w�}�v�6���xֿLVxT�p�BI�� �J�A�K]6VU�׻�6C�<-��jH!�oŹy���	sJ��k_�B �T��ݍ���� i���p�֎~�U�F9�S�sNz���1���p�3��V�O�Zٛ	E��&n	9K�佳'n6�h�0���f�_+C6�SK�ֵ����g��M�l����.���ew@{ы��ן�Dj��`Rx6�BQ��h W��}��N=�Ȇ+��d��5�h#>L�FV���/��g������<M�׈����l��)��p����~2��ү��rBD� ӴQ�:ELzjh��ه���t��c��њ��D��1u"N}8��:��K�\̱�`oA�@�I�`������nv�A�@��˗-e�!Ⱦ{�y�c��<��"��+�Q�[2���H�KP.�UҚШu��TRf��duw�	�e�����"r$V���7;)��ΔvdBNU�n�{+w˟5���[IG]�(UO}Vrf�3rK�EC�4$����Q�`wQA�~� =v�1rw�iC?8��^k��2~�]E8��8BK��ĥ �@�x�gj�7���¾m��b��_���τD�8Bs	���/�DY.Zǀ��zbFS�>%�Xf?��8�$V"�E�(T���ZH�b����{r��E`i<U�iv27F�������*y��"7_)�G�ĕ� �HL��=4oB��av-(�����KQ�<���saLU*U� �硸���9�j"3S
�n��;��%�K#����;�����������&�^��"��3
]��Uy�`yL�-��o����Uhn��6�K�g;Z�6Ʉ�5�x��K�4j	ةhx�sh�	@ᛥ?����#���*C��a��f~����-D��֍1�e8�8��_��0h-�s}�|'�Y\ڐ����~7Y�=y�����v��H,�I��@d=�.h���.�ւ����[M	�~>kV5
��+{�*�X�q��^7d���"��rg�xV�uRh#�l�dF�u�AU�xE�C�?�IN��:�p@�^����m���p�B���	�!)��`w�_��µY@	f1��g��}�Af���ȫ[+O*�Hz���'7��y���h��+��Vu�^'�~�)ދM��3Y)�����z|���-�7oH����RF�K�������A������N�֧ؐ��6�h͛L �˓��N>#��!���ĭ���-�
Iiw��׆&��@���؋�DA�	�\���f����A"l�|�܉�����8��T�W�R�.�n���{���􎲝��[�V8��������NK{R�943�����n6��������B���m_ݦ�n:C��v�rZ�C*�@��^��x���SZ�c6(;������m�$�'g�� �������^�捅R�<L(8� �+b��<^#+�w��u���V�������'��)�B����%��E��V �.V&8�d�F� m��L(L�]sүO%��T�B��������~�A��lpDb%�dnh2���П��Sj��T�������E��P�\�H�w�)OO���Z�,�R�š	��{)ܳٶb���@�60�@ĦR�$�P�"auYU�|,�ٌ�4m����8l��0� �_p��|�_>Yۈ*#7@�S��{��I�Z��#�8žmc�
�����2�
�5,�V �-z����2;��l(�}����o����%��ׂ���i�����X!�ʟP��e�=���s�:��V��H"������j/g���mG��%�ᦝ�?�$Y���¦�V���D����\**�5�+��ðWP�^'��2y�o�>O���f����\���>J���3A��s�PP�TLv�U�[=���J+u����<��?P��(���T�h�N�f��T�)��Nh�`Uj�k>M��?wT,��b��NS~7�dj�/�H����r2+(�)u_7�����t�����O�X�*'l-�M�5tUtG�.w��n�����6_M
�m�3$+��qfS��U�^{��2w��u(Z��/�Y��W��2i�8Z\־Ό�D�㯵���z�`J<��g%7�
2&�AF �Wik�C��"��T�˚���"n|Z9�)\�Hej���fǍy�ɫ��:-gc�/Ώc��n�e��y{���ìCV�9��M�� ����[�,u�Rm��@��K��2��	��d@zU�<r�t�៳ /+�l�)��ْ��3^����?�������p����lN���sƞO|m���ɕaQ�>_q��#���R���2.�bf���M�kPy�
��i���\�p+�ٌu)ٛa4�x�t�@Ìݕ^�
% /�~>Ό��.l
F��hW���xT5�;H)�]�ٺ(��鈍��Q��d}�:��rl\<����?���m��@Y�lɧj��ʘ]]~\�~�� /�Y�r��)O,'��q��L'�e�v�LG=Vj�Wd�b�b��E��&bĹm��d�NT#���_�v4<V�I��QCY���!?�����:�W6��x5^,�d:ZMR��\���bY�``�������^�M��{�K���&����}B&�8J,��-����U_����Tg��G��X�/��
�N���q��6��rQ�ش	�݀s@*ɕV:�Qi(�\��^{j���Jqs:U�,Xt#��,ZZП�R���C�J3J�'Ō�د����+O��v%� S�v*-�¦�ez��Q�&��&�}}(V/�2��ؐ���=/���<o�i��.Mܢ������o�Ein���#Si�Xީ`[�'�.B�����?���&'D'�АIz5e�6����~�0vXN�Uo�`w�8p�k�L�WkYyЬf	:���Y�񫹋�ORG�}u���S��4��r <��g$��#�[�؝Q�=�&sV���I���]����6�su��MXY����Beu�D������yF��M���RS��R�C�'��eXγ	85������#L��#h}�ʥ0K�!��-��4H���,�@,�7v����bJS�Ґ�!���<}���H��G�x�'K�L΀�}�#�������({��Sx@0Ӝ'Zg�}��=}�CYL;�	�W�) Ei���`��,�Mw���(Q��hZ�Oe�E�7�\T��[�EH�|hHQ��|��Aл'�|��D�JJ�ȸNp�ֲyU�Jd?��shw��U�$�ы���K�Q�{ �gN(D\�����r@�[Y�4�KM!�Ě�0�?#CU��E
��a��̺vEy'�sI���*]iu5���1 �P�ҡُ'IF/���:${�(dR�ϱ�V�ۥ��Z.��>W��������ψ���2���Y���0�=QAG�:��=G�G��p8q�M�hQ����U!��X����O�t��HL� 1�y�Ͽ��x�y>ux�K�f<����6x��=|���㻑w�ޙF�;uL�*)���˔|��xi�V<�}tJ�(��ܗ��JvD���{��%�EF�>�Z6��ѽѮ(��+D�m���8���H��#���{�ys}uoK�K���C���9t��6>'�t����YH���� ��,�I��9ug[��銰�D��+�؃�5�k�	�O�ϔ��q�O�-�ݘ�413��N���M0�r��9�̻���q�@�O֟�B�{^�8�>^��b����s���YFc���)�R��^Uc��f�,|�">��j��ٚJB�d��Y�#q���o�ڻ[悟��b#�6ӟi�Y)t��3�D@�۔��]�7>icN��-/������!�P���C�Ω:y?AT4MK�i�#�,-vp,y�bа7D��{���N��I|�V+�i���p���h�l��rX���#�π�7�rL΍�#��#����mH�QmJXjqa�E����pr3�u?�¹yB�.9;Tؒ�ͮ�>���?��*X�����a�	FX�+��7eӾ���8z���^�˸ꎄ�^KUpY�5>�_���ɒ:��)������M-Oŷ(<j�\f��u�ؚ$���	��������Fv��t�ֻ�v[�Ŋ�t�}�g�k��FcdSo����(xs&�hH~h24��0��P�=Ӫ����\t�>/��4SD�Eѐ��Q����'ɘ�+$|���7�"N�0~Mq̸�s�`Ս�)q�s9T�4\����G�/��'�)�5
H��a5e�ck ���,�뜫A��q����v���s���������iĸ�-��YQp8&�hs!ؚ�&�G�����L;�6ݎ���w���M��<PCa�K,=[X�bA�N�wkvGIi���a�u]���<�v��ނL_>o���o=�מ��Џ��wvu��V`�H��"OT��[#³Ӝ���cō���u<"�����0*aT���kv�?N�z�o�F�tϽr����	��o����}���|(��������ߣ�=����xxOQ�U�؉qSIgq&��PK�u�7p���|����a��Yͯ׬@�^Ab��l�8�U9�~����<e�8�D��9�] R���x�r��	�n��� ܵWgg��IcA���UF����E+%Թ\ۂ4��҇���I����#+зL�)3�{2rO�ݧ��V��P&<�+�E������T�9yѽ�OpA���l�t�3-*�Os]�WZu�����ɶ�X":^)��
�خ�Tݢ��s�7�_b���'EI1��� j��0N�'����`_|���Máw�1�Ŝq��Tŏ�=�@s�L��c�Ɍ�k����4�k�:��1�/�R��KS�t��r=�jnmS'�~�Yd��QZ��T�������pq�)	w���:�X \��U�T�D!��h��q8$�>H�T�`Z?��x� �2���¡���)�;3�>%h[8w�#Ǽ�X�\��)�P�pT�5й�B����^�%�o�
G-׌��z�/���r���'9�>��RE`,��}z�R��|�r=����}�qmI8ʅ����N����o�}�Q�_=ɣ5�4���E�������;����9k�xkI���b����;�k�Vh\�)�M�Sس��ǈt�`�ϛ�=���n5����s�9S��K�RfzE��E�"2e����x�l��"p~c���!0:�λ���7�.������j�j,���åw���

#��!�/���y���c=�=�-K��|#W7�~;)��M|�<�3%�{�t7_�m4����4�鎣����:m$w}�����?���ޥ4<M:��i-[h�n�5�IC�*M��2�
*�X_�w�̤R;�.uKܟ7qPk�RVfh�zZ�<y�7�IM�����;,�E)��s�hhp�C5�Fp��G>�ldnp��Z�UW\+5�>4��c�u�A��k߰�W�Q��3U^��p�/?5m�S��t�5k���h �~�&����e2"`h[�Π@�3Ur"D�k[0�F���"8O����E>]!�İI�@pƶ�/�*��H��L�@��E����%��!%F����*��+�E����AQ�V�@;�/�	{!�8��@�� ny�5��$����&48Ǌ5f��)�H�ڂ��J�YɁf�(�'�tla0Wkd?�����AwnC�g��9r� E.�S��<Y�qm�W�ɆoW��PJ������ɡ/Q`ze ΠJPb�"^�B��e�w�5�ۨ��=�i��ߵ��Td�U��c�?'|��/n�EM��,|��P~8�ܼqPA��(���&�d�춮.�_� 4W�s���:�y���3���SU��F� W��(%Q&j��QA��S�b���)13ɕ��Z�*��r����m��p_o�l3i��kmo͎�]v��$����=P�41��u(��S��ދ$68��	_B�@�	���`�7.���ٲ�5<&dWq�t}\ v�}Q!)��ҡ�AفT@�E1�Nߍm��k�@K9�_��phz��� h����}�5�L�	k]S��b�f4�����7Z���h��{�m�W���=G����Wu�m�������Se�@_��qǯ�}�Y���M�2U�gx:�k*)�)�\k��F��k���¡��i��5n3��6(I����n-_"���̊[�P'�����ʩ��(/���Q��Gf����J����_�����F9
�7h���iE��m�a����?��!�`����t���+������� ���cb���,+��C��"�鍋{pzO�M�U��L�c
7����n�B6��g�f�FID������E˱�&�?�Y5���2��&3&P�-��_����	La��2E"���B�@�Õ�����I\���7�W���L����cvC�V��^�x���Y���)�L��G"��ϾU�����!�D�b�eOs�d�<rG�q��Ak�fV���$t�ۚ�A��;�2>��d��@�7!����'�|��v�0����w�Xp�4 R���?GZP�征]|�?@�9[r��$��w��u��[
��q��pQ��1����~�V4D��+���M
��j�ٶ�l�0 gV���ּ�haa(��y1^1lI�9M;��7t���wK������ ,����R�+U�F�!��1X#�t��QX7M�+$���4��r=�|�:���֩27�c%�$��#4���i�F�C�Y$����8�g���9�3!酆�LԲE�DH���+�RY�b!k��H����Sv1?�=b�5#
�ˁ��,�g)��4M[�cE���k������Y����}0���ku��3,в+�j�xE���%r�0?���(ľ���ρ��C�}�T�{��H!�r���<��������n��{ql�p�iETpK.�BY��6��M�ov?�g���,}��K�\�������r��Z���vW�����b+����Ј �A_s����pZΞZ)>ёzM����r�I\��LpSga1�}���b�Ve�G����4}2߸�UX�0����-�w�����]���M(0Ǳ ܐ@LꮊQ3�x��d�tT~�l�=ֿ��a� Y$.�����V&����E� � �0�� �?�<����ЬK�̙��^)��((��4<��ώ�^R�E�e�+�p�����-=`:�R(z�;����3D'�9HjEE�< s���k��V�e��H�H�ڋA�T@u�vi>l��M?L�b��|�٤�I�ј#C�|���sV���"$䰟 f��iZ��g/���,R]\>Hf��H�I�nX��W��<�
֨�:����$����C,�η�-��RTk�8��j|�]��B�B��wk��7wV �N��͠��?�	�V���7F�f�#�ל�M� �p��DG�j�F*�o�yp+t��6[����Kw���k1��]Y��R�/��~Tl��S����j%�k�`��������:"��f�*~�h^�Lg���s`SVp�ۻ.�	��]��&���D��5���?�\=im����a�����ؓ�s��1����u�h	���k&�uMĵ֦������Y��נ�J�=<��	�<��Qz��W��ȞN��ZL�������ۮ$�J�x*)����h�W�T�U�_j�������Af����T�,V�	�l;����&o�фoA��$�����BO=y�����	���+�U�W�~�!�4�R� ��s�U��zx�>nt@z���.�z����!��y�$ �g�F��dme?�Z>��n���tC����s`���\P����ɰ �<!&�8�J�}��_�ll(�~Ɩ��_�G�m�A��{�&��2�#$,#��n��b�O���Pʠ�譗	��*	Yv;�LI�(�����s!�Dl��=�W=��$x;���X!�4���9�v4e��1v�7#�%]8�	�7������ TU)A{�WQ^���}�.C���
��Z���r_�/�?�{�wj]�e+b�g6���D4u8��	V�u�(6O��ʷiLl�7Mo?�F�S��"Gߞ�*5�����n�ϷK��5�5D���P�6Q��,�/	�y�	��%��t���/i<��+#���&�G�]�/q�L���Bc�K̇\O����DV�����e���j|��0Fj��{���9���⌂n[����s�	���b���)d���BK�R���˯CkP�!�p#@Jb
p�o�g�=����b���u素53O�3zϽ���@_$)��O=��7sm4�*!֢�$��s���-�L{%���z@�Ř����*c�:�歭�{GGHiM{K+�� Z���Ĥ�	-୓q''�;Ej� hߢ��y