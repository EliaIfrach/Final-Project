��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
�bR�{���t����^���%�T�9�;2��#�d���R[i�h�����Kk`hp�襍�j��������k�e���w7Ӛ���a=��l���d�i�!-b�_j�G��	�!9�ݫp���7/��?% �u����td�㬷B��Xzz~5���4����h�C��mȪY�������6�i,�OO5�ct���
f�$�	2���>4��j�պ�yQ��p}�F��,�(���$n��c<����8!�T\6a��ŗ�=c���٭�Z;q��8{	ʖ�w"; \�W}g ��Vv���+0^!�N��x������Æ���΁�L>�g�Ŗ��j�sSY��i��9��kƀ���;o<���^%7�N72 �]���&�z!������H�h�5rD(���JU�����˞�m�DB}��1�O����j����ruxBE�6�O�
v ��y���mȇ��!QҔͽ��ʐ]я��u�5~ġ�����qybs�Vh����Y�O�G|�봆G&3�BU겊ǫ-�&Z�Yc�:���f�z/Ѝ��$��7�p�:��\�1����̻��@�%7,j��B�@B��Cp�b��O��_xs2ymV�� ?�y	X)��S3:ѳ���!����G�V���h��[ȃ�@:|�O����&���+����;�־d0��P�O8.W��ԋ��ï=3���<r����Q��a���/ˤ^���?��6������y�k䷸b�
7�V�铮�����N�+�hZ�J�F6�<Èw����8'�R2$Aa����b����4@��q`m?�mz� ?sA_N�nƅ�{as�H5q�z��"��'����$�z:�%�E�ڦSb�+��Q���`�}��fsj�d�|�2��Q�����5fzE��i�,����VK���f�D���:����Z?ɀ��$5���~��K�����(��[9ݗ��!��{^o$�a���Ĭ���b�S?�!�q�?U���QN���/�\U۹_>�*�A�>��Q��F�O��"6������ۤ��/��6�A f�D�����`֤dYd�/��U#���+�PS��3H�z�+R�Q��e�����M��ba����	3n�efL��W�({���Aٹ#u�B&W���:ޱ)�L��q�@| 
�bHn=��叝�-:�/��g�Ĩ"��p��W2�pz)I��}��{���Fڸ�BU6�@hY��p
g�����2AA']���O$�k���k�(�-�x��ÀLp����x"��ϣ��Z,��(�l@܌��*^�C����ɤH1���2Wp*;��w�㢧���&���%��R�'�t�U�G�E��!��e����LԪ!��e�e�T�rIخ"Yw�kƢĴ�X(����x���y�ܼ�
��)��w0�-X����#:&VЭ�hG�����	�nW����.�P-�~���M*�R����}�i �[�b�p�p���M� ���j�(����	B=�M�,{������i|I�ƅ�KU�`j���֢�ھ_s�����+$���I�l�Z���;�� C�7V�0ǅ����a�Ӵ�¶��׿'7��V��@�xvWir^�?�S��3��)���Wo�a�QmUTO|�|0|���k�]�[��
F?�jث��M���HJD�8|4-��U��i$������?D�0������#e��[��4�i�����3i�4�9-��-�潕�=1�FRE��7��?
�S��;�����J	h�T\�Gf�B�E ����#��C��<8��]GSy[=���*@�p�����E�bU��� ױ>�I��y8�r�PHg�W+\�߀c��P�N���Q&�f4���7�� ~n�'Azi����a�<��e��A`�@�X8�s���=[�#�caBXpp	�hr������t�9f�.��dcg���}¯V�)
c�\�wF3�?
�U�N��I�}־�
��h�f�B��${�.��YȲ�L��?,l&��=,�������U3g�i��M�DڰK#��!�ܡd�=Y�s���`P����Q�0�_�?V潠H� ��#���Zd�p�����f'�g���J>�p
���{�ر����ʍ�M�MQa���p�~g���cO��Z������0��q�E"�
���̊�� `�������r*��������]��(�(�c�#�d@�(�р}���؃u/��b9fTNw%,�`�� �q���9�>��-0J}L�P5�Yۤk�Г%f�=�0��@{2��� jT�����zTH<[!�����{��~p���J���1mU��즫�iV��
`�N�7�,č>���]�@���u�P�>���:f7ўA���q���ճ�o�-�M��E[)&��Sm;�Jݫ� ��}yqK9���J�W��P�̶W�zltu�w�X�5r죋�4ޣnh�M��B�6\ұ�3Nk�3��/���C݄}!��an$�!H0N˂�0����->��V%�R�v��v�`$l�S���K#���=.��C!���u�w�\^��B�^�GGr$uLsQ�7��W���{.h�D����K`@�b��ni8���Y����	�m�cMk�Ow��H6z�8��.;�������^�	��|)���{�Q�.�-	�M�8-*���l�'%�Ŕb�b�c�T�#����e#�d�G"�r��)�����dt��'�����^ڬ`y'��o��`�(��O��T���Y�ҽ��g����;tn*�E#�I\���\� �n�N�͓��U�����@�fb/o\j#ؕ_�s	u��e��jp�u����@����ɝq�L��[(�WOh�a���	�`;x�<�0���辀�I�Q�4Z'��cr|��]5Xy��~A��Z�nU[��*k#Y1�W�U)ﶇۤ�L�4�b�k����/�� t�n|Q�� �;$e�m��SF+��(�`d�Y�����Qp�~���,�<l�̴��bW?Ij�A��z
9W!��+C,�Wg���Dx��:I�Yeq :ɚBiAIp��KY1�-�~Mԭ&��l����(�����w��d-$(��g=����g"��R��s�I)��p��zZ ��mN5�|�� ��OQ0bT� �/��ɄH^�����zrm#����r�x������@H+� �HT��&o��xR����w��JY.J�R��8��k>^L�"�9�2I�G-��H��Az%]*�U�k�{E���.��d#|[C���pfB�e��B;X2����>E�0��ܰ0ATqO��M.l�#tv��<�X\T����4Oݩ9��'�ӎc�C�����-џ/E�;H;�$K����Ūb�>�_o�89e���<_ �'L����P^�� �� ��{@�$r���V>`��;���B>ő�l%/�/`]�4�Yg,�c�SE�~	�f����je��@��/�Y�<�m�[���D$��:�R���Ҍs|�'�=c�"X��
��O�����*�F��?H��un����"�n}�|�Q�4�܅�E���Er�s��h�J�2(=��g۽F�=3v�fg��l�*a\��65B��Ҝ�g�=n��/����6��=OW�X�}�0�9c]�{�����md��'�5���c�p��ʑ��7ꮬ�K�E�Ť�����2�3M���@	�@���DM�O�C��{\�~w�0a�|���/�X���"�����cq����-��S�c�{Y�����g.�g~R��� P�դbRF���5O<.���*��x�2��S��V��!bM?�,�[�&�Tps����W��tg�&42]���:�'bt�Dg�˷4���ځ�� �+C�Į����P�,��O�B��11�5.U��'�eYW�o>��:�ޕƑd3g���Fl� /w�a��e��Ӌ%�U��������jL��_�r���	>�Q�Y����j2X}͇7K�;T{�2`�2��	�Ɇ�>�[�v�>�eX}B���?(��ɺY�a&J����hy���G������=�b�(�H�g��P�b��
�,_��mcɲ,ۏ�Y�4Y�#?ٲ&Fi���~ݛ"�e�)R,c/�u9��ݮ�˾_{�`g�x�\R���g�U�c��?ߌ���V��ۛq�����z&7A=�hfHN�^g��vE�o�F*&���x�*^3`<A���a��97��z|����es���K<"�z��sq�K��P��DW!U ~��r�v��f��A�Z3]]�������`�|
�KG��c�o��5�|��ؘ&�ɸ$�:F��jy���_�Ty�d5�"} ��R�.h�?f�;F�NeL��͋��+;>�+����˗5M½����R����,��	D;�Q��_���>��z��$$�F��'9V��[@V]\��|L��\���Zx8kP�P]U��+e�� ռ�j��l��j&�I徤+��/`�`���.}盼>�t��kb-��Y�e����X��i��u�o�?2����@?C��D}N)�
^+M�nI�2�����#�/sb��Ȁ�DC̱��t%da�T��>j"_�b�'��q��+��Z��ӯbPZD��ƈ�D\ԥ���m������ fQj�P��L&Zd&W��p]���,}&$.c6@���A�o��~�>�hm�(���s�+5����L���I\\e�����n{�������'o+\��+�*�4�������3�<��ѡs=���	��\�ӗ��`�_���8���4�cߨ���i��y#b� uU���4ƥ��r�G��ex�W�sy�<���X7(�&�R��	�1�@R���U��5[2�*�� P��<f ���Y��)۲�/�2k��:�3�k��bL�\-� �&�,�~.�gs���!*,�!�����׼����{7���������p������rl!�G�V���5�~���]��2��#�'�SrK��R�J~�j��:�.��9��� ����B�4�� ��z�3#:ґ��/��m�X@C&靡�����H��3�������6�p��؂�$�4b�y�1F��[��E �T���i�;�}�u��!|�U���>s>�"�A���i�R�y}1Ʌ(�H����cC9�s6��r��u��Ҽ�Q=�(�M�!�r[&�|K��ڦ�/. �S=������HH�2�J�W=~GN��l IB�Er�K6��"�%>]�?<�7��	{Vi�95E��b G�xvf�]�_��-N��̝i(!m�x�*㈜yG�~�Gx�7�� ���im�FO-i�[ǹ�tae[y{B��u*S�M�z(�/p_cp��	�I��U���V#��l�^����d8�H�bh��i:���)xC���An\�u�lb�yO�m1�?�����1��&���j�ITw4��y���xq��g׬�����2���؝��=L1oXlP���б���Lƴ�@�c���5���Lj,#8��W�ۡ�q��٫�QY�� ��p\����5� ��8�Y������j覤LH�&#>'4��ѽ���5<(.4r�'<�@��ѷG��o��(`%Y���{!�hx�@�ug��ꤳy����4�D�����|ؠ�-�E���ҹ�i���Eχm�����M7����k��L�ٖag�/����.@~��d^慪�nC�Ut���b�<K���:1b�D0⹸�"�]XF&�� l:���İ٢�Ch� �6��,@�����(W�S�(�-D@�i23e��7`���5ǁ�G߷������?d̠�p� �#����y�,Z�.0��-"\+0F��i��	4��UN���)G�Z)`u��kZ���x�Q���E�c�eO���/f��cܞ���%��-FA!u�HӞU��%7��C�\��B��3��jG���V���;q�3��M����(h~�K�r���\<o(y��aj�x�o5������CH3b�U���<�`��W�6�`]��
����z�d������#���,x�[��G����l��jRJ���G��a�G�}�X]��e�^. T������d�jn鲗���.�!=P����K,�T�o���h�����
��Cu������ZDT�{�V����v��U`U�M�`�ǅJ�	�΁{��#��?��lnnWy)������f��S�#�A���*�L/Pp5��' zV��`���|�]>���ٲH���r��O��
�nP���8x���l���z'�,O���z��0���?ο�c������)V���퐦˹&���cs��o�RP�a�1^�oZ�*�˲�,A���\j�k������L
u-y`q2
�1]�8�9joəϷ��4����C��Z5�4͜�J�f�n��?'F�5���T�I��$z�����I �A:�q��T��ژ{�����4g�����2/w'f(�?��M0dg�^})ȱ�5��=p��,%�� �"���N���h�����C�i8�w��E��ƒ����Y�"�P*�a˃7c�7恐��������E@=1I��Z��U�'�Ƥ`dg�ه���0XX�q�,��[ ���.��p�3�W�s�W����m�<��0�����י[�@��]��d�����+�-{ح�G[֧޼1�A���{}W��c�u����v>]~��Ɋ7�� �ҁx�O��e�X�o�_�#���� ��zW?�؄���- �L�wu��Q���Z����%�^ԧ�����
E�;Tfﾤ���;��,��#� O����������ɷ2:�\f�(�4����ਲ਼�� �}��0,�k6�Q�+)��C�b,��tpmCeE�=L,	��T��cǉT�5������q}"�r�����د�ۼ��6��O��"���*�P�x (̌2k�&i�����0C�����H۰��0̋�ie�T	� �L�J�v�"ɇ�Q�~W���'p�<ay����Z��J���o�,{+X�r��-��[zx[��A9Փ���r<&Yz7?�vuE��Q5~D~�xB�ĕ��yJ�����}R ʠs�x��|ς�I�?���}^��H.�
	F�b�3`�[��&@�ifˮdet��9���-w6^�
1n4��Q�W^��Ȳo�N�>���t֟eE��e����R�],�E���p�T_3sIF'�J'���,-zNK/�_����P�J�$#�΍�5�fRka�WJ����%��M�� ����@���e���X�,{#!̫Q���j0�ݽj�L�����H>���>EO��Tb.7!����|�q��_������c�2�i�,�3]W�a�	�@�����4S�I�g�T⦧ZB�����Sj	j���w��a��	�-g�`�%�s�.CM�P�����OYF��߮n�8��?��gK�́�@�',7 ������>i ����(;��n��)��ͅ���T��3ZQ6��ŮF�d��>�����}*Ju�w�HsM�`̸����6�R=3�����`�¹�k�!*ޤJ�����Jsg��Xx�{Lj�A>��i�/W�ތ��_V���£J�k�-L '���pZ�@i���|I��_�o���ӽ&������!�Ʉ.�~)ξ�WԔbƫ/����*}��&�2�aW�fJ��(�������%�L<�s���.��q�NpaG��y�����^��	�D�o74pU�6)�B$�ٛ���N���땈�ͳhM�7I;?#ތ�/��1,f
�w�:����	y���h�,���Q�mQ���K�D�QBϹ�M{���^�6يvw㫠�m��;�����"��MR��9	����)���L�ٽ� :��Q6�9*��_�069�>�.���u��P���eA2.��a�z���5��{�?��Kv�Ŷ�h��>�}���<b;!�?T|��)d)Q�&Z�ڑ�٥���R�`m�.�H�4fo�'�ա��Q�;ǣ����L�FR���W(¿�=��%�y��^�P���JK@Խp��j8�v��4��[���C����H&�� �>����6����`b`z
Q|�M
��J�ѡj�AE^�i���$���i�i�X{�G��T����j7�@�a7h�-}Cv��.=�
�d�!z}s����c�Z���|h�ҎN��(�|/O��'CLV���r��J|��3N�M��8m<�2b��lu�	$�2�"�U�|u�u�ǁ>tƏ�!˔0k�m�3��,O3J	��ye�dPV�HN��)9��ys�����������BP�u�R�kƇ���i��r/>�e����F� �K�c�X�~�G^�G
��=@�ڻB�Qf��c��'��婟����9��"5#tC��񎐮�)H3i�l�ͻ	�"�7QeC./�ըҊ;`'i�oJ�8)���42֪��&�7t������4��E!*˻9!XQ� �z/^"�5�dS��(f1����${�A�\����]��m�zL!d�~x-J���^�m�T�����M3�-QtO��䰬X2A�����A|/Ɋ;���˘�E'H����,�T��;�k��|��1�´Qi��Y�]�՜���2��u$��H��-�d����V���&�~!��~�M�<�J�M����~������k2���_��7�6]��S�h�rm�fi-��h ����f�$�% jaR���:�q��7[j\q�)�ˆ�^zi��e#1� �W����/nMX� ���( *���0��%a��9���;��<�v�nM�?�N]�uƣ-]�QAW�n�J����F��/Q��|�6:
X�� V,ʰ��[.�H��.�~3�P��w3�9	�# ��d���%6f��c��Xy�]�:��T�J)�I�$�Ts��:�7�Ǻ=�>��˩d�	r2_����(G��< �>�fV��fB�P����*f�D<S��b
��3�Ҵ���qA����H�Fe�Y@wal�}����	3�D?�%{��}g��<��(��.��؜)��4�(�A�+��l����.C�e^�y|�L��K��[l�`ؙ��$n�~��Gb�P�z� =&��R�����~!�o�!r�|P8
}�:V5���zcdFq��������)�cGb��.�oh�3�ݭ$@r!�[��k�\��[�� �=5v&�:�`��91.�0u7��Y�침)`�u�s%�Ȱ)>^���m�eoе��|����_қY�KL�>�M55�pVn�����L=����1�c#-�g��2+��ʱǁ��+��	FQ;l����7�����H�V������O��w�M֣̂7Bx���ZC��O^w:�Q� �[=�����<Uf)�0n�,�P1���-�@U`��Nv�a�/�:y���02u�K�׷��z���q��c@���x�~�y)�!o���}��:J�ͳ�dn���V�G�K�I��.V��Y�m�����x����P�?֩���lP�$QXާYV6Т��k��X��vS�Kk��2��:��$��j@�J��y�Q���d�f�Peo���(���u4ƤP����m;�Zu@��JH� �m�'����m($[�"ݶ�^�W��?��H �-��	�#�-P}e|�95T�h���!7�&�j3�s����Q�W?�1KX�i�W��oL�22S����	5������q~l�w䛂�]���� hp������5����J4��M�W�v�h5�z�&v��]���c�A �0sDI��Ʀĳ�2�8�FV2��J�ӎ��E�B������%á�:��,[��`�o� 2EH:�E�z�u*҂r�1a�����c�2٤4���V���aky�+���t&�_R��qn�2�'�5վ�f����r|��xah1������q�G7J8���zt�S��;���{�P�/�wYV��D�6c�ۢm��>F��rt#��L�����%�F�nz_|���S�����w��*�q<������F#�'��\�j�{I��sl2�Nz�LP�d|�^����8����>ÃTۜd�,�[B�9=�|t��aC0qcj�@��gN���<o+���ڒ�i�J~a��l��+�N���'}�S��`#uZ��,�[�	.���o�uY�9��p��N��>��wEG>�E�[��P��ߑ�S���'�����D�sR95c��p�h7J�I��u�|V�uD��{@d���ߵ���2�-s&L�YYP ¯V�25�Qi,�.Q��ۃ�5��R�u+�l����f����8��k.2?+Ԧ��y����o>��ͼ�;�͌�c���M	g������k�!����Ԉ�i�l�������VBɜ���Z��_�NҨZ���Ε�J
���Pۧ�f��lh�lA���þ^��l;^�o|�KJgD�U�1�;���M���p���z�{��͍�p��qn�u�t�?~�pWZ�z�����8���w�M�R ��&�C���8鈣F m�W_����<���p0>U^2�ݔ��5� ^�HЮ�q1�U��h�������.Of�lP��D��v����޾6 r����cp8����P�m���"�F�\���uy�;VS'��:���ұVw�q���XO/��3U� �H���d1r�,���=�z�?�j�&���QD�h1�t�v];|�}|����ڦ��v�Q��i�K�:#2 ���S�(.�nk+����� ��7�/W��QϏ�~�_7'%l?�2t������I����o��Y�KT�9P�z%L��#�=��f�U�� _�����@�	"%1����ӣBW�����u���8yϿ�A_^|�_�^�##p���k����\q;�����W�o�KJ>��ʘ�L_C�2��q ۡ�A��0�R7�r����bi�1�ӌT���ی��\�˪���3���Y[��O?'��Cx5�\��'��X�RIr�=.DUU���£'S1�o�L�ݬ��}<�].V�b�Y��h��F�,�O�N�ڼ�k4���Q�ۻ�lX���\�ϦM��(�|Fd+�Y�%�����m3����ݩ�â�U^���&[�H �-����+'�haX�	1�D�׋���jҡ�~j�Pfciĥ���̢d�EYw��w��4]�8�R�3!eP��D����% �Q{Z!�{=8���B��a	���~�r*F�������t�H��-Jp»��ZXc�v��f�D��i� !{:��i����N&�����y�KT�d-c�hA��No�	��&z��Ť��
?Dia*b:�aW�Xi��M�g�>X�A���؞�W=9F�vs�anN�ځcO�r��\+0+}��D�1*!vSƊ	k)�w�z�8��<ر,��:�%_0'��?�cF[&���d��_�ƈ�E�	�½J��1���C8�y=�{�l���1��Ѳ��	�h�����u�3E@��>�0�ҼY���>H$x5{E8������rA~�?b/9E_r^�x:�i����o��")�⾃���lH�^���he;�`yC�{$	L���Ih��b%6�KU�*�#[YY��K�����gq	D��Nh�D=�98M�6�Z������sH�� ��r��ϙ��o��әV!n���7�8R3j��S�~x�A�?~گ�ESc�f啎������q�Ee�ӐdAX�L��OIB8����>T�<�_����	y��TZ�;��D������P
}����f���5s����
���6%�W/1VI:�s�>kn�	Z3�Yz¾�V��C�{��4?����R��J�|�vr_�:�]/���y~�c�/��}���˼h.NyZ���;���@���y'�o7��x��N�R�$P�l������H��I��
����Ҫ�d���h�a
��7�6�~oj
�،֬0>�¯D�=�q��Y�����D'@{N�<`�Y����Ƒ��1���?¼G�1J��� ;]���P�\���͕�V�'q��%�u�}mȱ+P�V$���xN8��&�V!ӱ\Ww'uiBj�\�o��[���\���@�tk4(����t��!���;��r��W��7p��]�p9y?诉@�J��BD֖0�ҫ�D5RQ����0(���mp������7��6��V�$L����A�<Z�y�#�4�QAo.QC�4��<��'7�A ��,��n�[Kr-�x���#z����CP�d�1=���A@�����g�M5�E�(����8%�/M��Ƌ���(�dB^����x�>�����f�N�d���?�.ڴd4���NVz�lk�"���>���A~ؑ>O΢kDH:0o�YJ!��:h��A�ϼ�����XG,(��8u����2�ʍP|slj��*�]{q�$��s��왎]V�-f�}>�*�4��y�M�ݺӖ���.��*|�K� :ш�|i�r�],�����udf�r�R�641W��f�hK�^
�_�{~�2�6�L(|Aa�H��	9�S������?��C�oe�++�%��1��ޭ��dȗux�z溲�c=�� O�Ԏ��3⨝�0z0�	W�n��Ж�*/z��w5A®�kG(���5M:�$Pd����m��/�ڧ�|L�C���յe0��{�:\�Dᡐ_�G�9;%U���V�$5�g�������%>�[đ���j���^c�q�<�v�{�}�Q@ɞΒ�����j�&P����OQ�"�h�adȩO���6s�?"4�0�1x_�j*��]R�Hy"�x�ҍl���F̩�9V�ǡ���3~���/;"BB�X��׽U�K��v4A����b;�M�Ck�Od�������]o+�󷉟�.ه(�8��绫	V}L�]25$�6�������퀿G�� ��h�N����X�_%�ۯ�k��fE	����0{aV�˥�5~�G:��&����ާ �	�s�z-쩢���a
��f���O�*��1��T�l]==G��<):Ȱ��)�,�����U��ޕ�M��&�gڧ�sR>��7k9Q�D��R,�]̹r�l�B��b�K����?N�9��.�E�Bʾf$4�(;���,f\�Gt�^��(:ŀ �w��̑�;�#�8������h��3�ھx	z�rO��	<��pT]�b�AH�F�GL�P����[`����M866��>J+{����u�I p�.0#��L�x�A�.���@T:wu�q�EB�6ށ�H%Y�I��dU�e�D1~��gp�m��͚�S?~��]qp���đ�׺�(�LE�Y'&�S�E8y�1��f��hbH�t{�h�Hz[^��t�>y��O�r�O�(6^��c�D�ɫ=hP�,몼�w���t��k�������~o���l��ɳy!/�ʺ�<�]!)��m	����x�ӽI����DZؾ���[˦�s)�Ò��@DKp��p��)�+٣���>Ƴc�oQ�bvx��Vf�0�Q<���S����O�-��My+G��]��pVGLܶL��v� Oz��DW��ҭ�(�o~u�T�^��2"�@f#�l��l�����/aⲨ����%z�yʐw�B�����/�����X���9�V��#PC���0lR�	��y��>����p�Ln�-��\1R]��֏ ];���4���Ⱥ�����ߺF�����%���Hw�A�)�c�0\�@X�x54��N�=��{c��e���:��)���}q*'�U�O{l	�VD���R�gQ>��!r���9c���tk	�dp�a&��X	� ���Ѝ۬R�0G�,1;�2�� ���_�g��B�TE��nϔ��v���s������ә��Z�o�G�u�s7f��Pǻ浬� ��^T�b�F�D�P��w��a6c�������Вh���$�u������wѾdl�H��݉Ws���_��V���9�ȱ3M�ӕ�e�=�C���l>+��=@?�e*��=٪�|�1��+-��a�;�tҿ҇���C�[ ���A�w(]xM�����Ԁ��y�;�����p��P�/��N��e2em�T��v�+!/)�9�sa���*=�����������?o�%��Eo�`��Uw��-�YS�j��f��y����I���'���?�.a�g�W�6��V����}ٜ�@�3�X�����d�.��諠��^,d9��Pb���>�G2ğ�������d�.��Q�0�I_I��~�M)@~@�ǅ�U�*�N���-I]Pd�* ����:��>d����6�M~Th(��֪..6y���,�OC_]�3�������5�Uޔ���g�K�aO�|��_� ��D6�A��݈Z�"����C���K�y���}��TB���ou���Z!�\(�I5Ԁ�p{Ƙ���l�A�DZ�Lة7I&��_�ֿx����ƅ����_w/˦SG���kHݤR���,SK}���2�0E\%��a�&x���{dA��d��L��i����kǄ�Ѡv�*�o9�:��:�9M����_��c�Et�z���l�%״���r���P�y�j!�2�˦�>�T5�<��R��L�/0"՘��P��g:"^��o<�QI�
q�k���B�I�Ս��;q��"�RSW��H�������o��{��_�Lb9�X�4��k�D,�}�A�3�!c�1�zP.R�'g�x;z���%������_���X��%���[.�F �+Ɲ�nH�/;�]|�	D�1^���{�8�(
%F���o�K����e~�:3�3��I����\���-<����M����\��&�	R
!~�a��IB�M=�C�CRQ�T�g6f��	X�E�r�?(��$�G����OOc�k�ph�L�iY�U�O�g��mǊ��a���X�CjӒ<QF�7��4?6:T��2��1,s��X��a�J�2ՙF6���t�R��-f����H��:��yZ"�-і6��1�K��^__8�~*86�O�ǃ�cU��KJ���i�[�k^�"�ؚ]D���=���Qقm�&S�����p��x�T c���s��4��-T^������C\=� "�E�Ė	j�Aų�����n��,�L#�ٗ�g}��A��j�h%�5çҊ:-
����Mk8��9B��7C�bm�<���<8^��|��Œ���=q�0��"��r~�-u|��%Z���&�L{o�;/N��x��E�x]�3�q��{u������p�N͓I�?|]J8��˒��% �;�=�)��k�3Bn��ul묪���5]P/����^/\q���Kg�_W�~ZU���>�[����� ̇��00ǵ�zz������<` ��%:��`ۃ�B�r4O���_��Yؒ�ɜf~L�O���܋x����q���S��X5\}�_\Ȩ��נ�U�3t�*�.M#�9J��*��N�D�!�;d_�X�����z�k����ڠQ4ع�Y�%`~�-��Vd7�()��hxӰ�c����|����?�l�"���<Y# 'a��H��@�����v�q=/��Y���ȑu�A/r�h(����q��o'�̞�S4���7�I�`��舩yWE�e�q�B����L�q{y��P�oz��GG�ѡQcv�F6rq��iH2�W����?��5�7o�o(�T�F�Ӑ��xO|	��PJ���u/HY�1e~���ܽk��7��G��v�\�&�4�6A��mEl]�k1�M�^>��U��iX\-�ܜ���n�3�#΁uĶd���
�yi
��P0b���d�O	�9�z<y2�IV!>�#W���Y�l�VE'���K?>&�㬆�8�
Nu�eM�N�dY�+;�F�B}�A]ɹ�[�HI��Y��J�qM3�w���M4�4OG̞W�Fi��݀v�����M�/o�?V�=}�ԟ-��ףI�\]]���j�����Cj,��cP0r��)_ˮ�_��Yuy��i�i(�N���F�ea*T��gU�V��v��6;T�!���^%��bM��.�T$�ߟ
�>-��᝙�B���e�v��Oe�h#/b���n�۝��Wx;��h�U�Cָ�TX4�.09�����7�rX٤�0�ȿ5j��#�lM��Tb�N�[��1]M����+9�^�Cr��a�%�"@C������"�T�Q���l�$tΌj�S�L�8�;��
V����2�	(̺{�z��(5s��a^��U�;W�,�ڢ懚���|  ��8%Il'8�b������4�3�q5�Vf��A4Cf�Ap4}�Ӄ7���r�rTQû��<bǁ���ɦ�����X�����0-�[�]�&�g�D���zp�1�hNlFK�������F��W�{sj�F6Hϖ�|��_��lE^Mӎ*���L�J���~���dP�oJ,D�����p�gKa�T�1��k�l ����o��k&KK)��'������d<G桥�e6�h���%�!B�j+&�E�4*���yQ���o�:f���D���G7k٤Z�_@���'�1"k�D|��ھ�g̛�U�?Z�<�A�ɋmN��D\���S������}��{TnO����s��M�H��p&R���usvzJ�����|�L�Dx�rO0�s��P�����R��v��E�[���r9&d�	cU]�L�}TE8�;ͮN!�x�Ϥc6�bE�ٝ&����Dv��/�?�U�ұW��%��z-�YF��*^��biᄋy�Eb�t"a�E�	 ��Y���L�E�$�VZ�VR�����S�3�|�4"g��
�B2���DZ7��ĭ ��5vԻ~w��ц����e�zp����/�m��̄T����̃��#��r����s JAj��/�y]0�}�}�i��b-����"~��>��lc���Y�U�4����&Y���J��O/�u\��
�(ǁ�͊�^� 5����w�I^�7o�N�J�H����hԥ503�(����)%������]J�����w5{�v�'�묤,]M=�R�V�cھl�t�2c�������cZ�׵��Z��&�
r��2��g���n���@.�����-��ݣ=Q����0��.�q�G��,��~-�N�	-1G���=�v���!�RZ��#�Q�%F� �C�������OnJ�H�q��3C�1˓zD-C&5�{i4I'gû���f�^ b)�0�.�x��+1��c�!E��� {V�ٽ+��Kٷ~ܩ���a=�屮!����/�e���T�\_fbt�n��rl7��6񱲦jH9�==fN���D�>e�>qQ1�ZAr�Y������b��P�KE,3���cA:�:��<�D4�ثWI����SE�F��;i�����NH�}i3P�ʛ� ����d��[��~q���h�"7����_rz\}��oK�euP.��@d���������-y��|�����	|.>;K��S�Lf�0��1�"I!.n��Ά�:~�`���Jg���חo��m�:�&@r�Ϻ��<�H��i�(f�T�W	��S�*3qۤFԏ��_��RZ�
♯zXF�O��x5C�%^��e�)�}Y��'��"���6G�I8T�_�����q�m�H:��6��j�%��d��9Н�gU2v}=�a�����AgqQ���n3�
Ǣ&	0����sL��
�pY`�+Ack��4`��{��7�~�zh��T�ǵ?֯ 8���vi&>������BG��M�Y}[��z�����^��n<������e�ȓ(c0�J�}��������+)��U^�#�B�g�酶֋:%}��Wr0Ɗ�X��w��	l�ҹk� ��1ɪ����}�}U�����w��+�æ7D�� lY�T����ņ�r����)1�B�	�p���͘ V)��2Cs�hڹ��ڭ������@A�Bd�m��J<�2�q��s���Z�H�9ml7�3X&�'�Ǝ�Γ#w��7﮽va��")?�{*
aG��~��d�_5@bW�ϴ��]\��ЃA�-}Tw4�)u��3� �8˅���p�;��HF��3l�-�=�ӷȉ�"�%p<|k����a�CE��׌�8�%�6�YO	��O���fp{� q}�D�c\F�	;!�)=CMBI�Y
/7=$�4W�"�Պ8iQ�pt<��<�V$�ވ�'����p�����"��VgA]�Ɋ�Y�� ��AF�-�\���#��->$�O���D��ԱSe!5�Q`(����4�̧�(��$j�mm��z)�qDe �w��4���3�����׷@0cS�O-}O�j-:t�^}��Y��,R�a_�BP"�
p�) �|a�S7S�g��|�uq®�Ӯ��k ��sh�%R������<D�[����u�9���H�X�)=jz2B��u�f�
�3��w!iw����T�
�3[ϰB���\u�1�Z�7�]�0WyV����>z��oe�W�SOL��j6�h c�\�ĳ��䲨�w�"�2��$�tF�YD*��(��44s��,B�ޯb�V��EҩD�k>�d�i�����~���.�q8��Á�����7��H<E�ɇ�,��:��]]��Dӱ���ou�Y��vr�CgZLJ���	5_i��g�7?è������S�=�����@U����Q�	dE)������	֏P�Ց]T��v����X���A饺��h5��N9�^�JKo��r�7_�Nz��Hj�/�� ��e��$s]�,��^b)骨ݬb�)��Y�Iނ�G��S�~s�WI��f�S�q֟n�s�q�ů�-�XzΊoK��E��W�n=��BS����[!zS������6�̞�SO4���<��P`Z�B�߱Et��7s�f�R�-�נ���7����$�-��0�Y�)?zP0�N�e.I�M%$y7+)��O��p1�ZJ�B�H_7p)W��k{(�e�T�7��f5,���\;�C�$�U�w���}���RI�sQ+�_��}'ctv�w��E�U2�-��-��o�tL90���� Z�#��t��pNKvk���^�|AAm9ȋ�ړ�i������\�g�j���"�aB�������ԭ0����g�z+	W9uߡD\������ �ͧFQ�$�օs2	��aȏ[B1djJ�i9��Dӱ���,���&���8�P9�@,��Rw:H�I�p�5��.�2�m�wƣ
���)�5�v�d ��g���dO�e�u���V)^Tg�?��|
�M�ֳ��0����jLr$Bc�H�{'�f�V�~��Ǧ#�u	��(-`��4�%�ݠ��~�	o���1��ٲ^�x�x_(/io�i_W�H?�j0bbY���Ǉ`�y<�xi����~_,�lo����ў|(�ڐ��s)�IW�}��bDV+(� |�JF�<��y�Է��©���]e<�5��0�=�X/�O#�0�5|2�����Y�dw��@�e|]Ǐ��[Pr��y��$1j�jo�#Ԥ&Y�O�#��ay�Q.v�u`p�T!Hk �!V�-]�#(�ίX��H�E֬�Yq��U���0���	ڂ����*H��q4f{qG>A���9^�D�܉�������V�s�رz&Z�!�Cd6��g�᰾H(}�-��t�mc�7[ �P�xg��<�$�T����B<v�1��C��I����Δ��I|ՋS�n��=P��AQ�Uu.��'j�*�:��b�����iw^r�a�DmA�N���X�K��xcXҬo(>�.��Qe�x*�O.dj�i�F��&��`;h�6������)kP�p]^�*U�
��.�9o��'�	^��1g<���_g��L��������PM�<�)�E�E3+�6f�����`o������x��V�o����U��e�K^�2���+������Ag�vM�5���4$jԝ#:\оl 9b���6�:��<�Ӳ��w���0Z�X���)T��睉�1A��f�?�S"���B1�qy����Y��}�ed�&�l�
J����>p��A�j8}�5��5��h��$����%��<~��a���՞Z��`��ј�ĳ�B�J��NY<�F��?�"�Ļ�t����nu�r�C:F���������"��2'Ю�e�^��f�F�˰ק���p������ M�	��(�My�X<Wc���xW��Sk������˶�P��K��oc_l�ip��;���Ck$b�Q�]��!�q��LZT������O8�`
|Fj�,��?_��'Q�T��N��&����${'���Pk�[�IH�BB�>��u>|��ʹ��岪��5����m7�<%L�C'�פ�s�3��v��Xк��<���M[?�iO�h("�Q��u�qH�a�n�	��I�l�o�wo[#��E�T`�셌f��Q��\����O {���n	`�~�z�$C�Iλ��dfު�-9?�Q�ƞ��8pHR$�P�$�3F��#�XY��@M�FB�ډ��CCĢM�G������v���Ra ����{K�Kz�l�^蛈0�6r^#ި�)��'�k�ú����+o�{�8����G��:���:�3�f ���&YtƬ!�`��B�q��E�}��H�]�}$�P�f/�0�Q�U����C�5�=-��$��U5���h+*>\E/�X�����O.X|YZ-$,߿�+�Of��d+��\���H�˿���t�� ��3�pA�K���1�%A�@���*{���icy�H��X0]{H\XVS�GU3M�{"����a ����TPY�~ ��<�1,S%s�$hZ$7��GD�<�k�A]=}d�ͅ9כ´���y��4Rva���Nۤdv�sB�n����o��?�z�y; ���cS9(#�ߤh��o�mu��DtpKR�}#bx��K��mO_�CK�op2g`L�A��kF�X�M��A���4�����s,��h�{м��{���$~oz2v�����ʐ3��i��w8;��m��A@L}��_�.2wWR��+8L�
�e������MA�F�� ��7�8_�@x=�b�\���Ǖ��<7�٣��� v�^Z%Ff�?����۴�-h�pBnx���{0q�r	{U�kGx�M&�XYf��qjf���j�UEfs�vt	�/����[ga������0H���d����?�j�n�2$Q��J�|�͈3���4��^��	B@^t�����ZB��h�=�k��i�Җl�#�=�է��B�0�E�j`������	n�	V�qK?g��]`+�U�#�]�@��1����:����1+&����Pr�ʌ�e�L����xڂ�4��	8 �0q�q�����N�~�j�~rk�ai"��
^^�fAx��h�q��E�H5`s��É�JR۶�u"���E�r�3E��p20`e��o��̝N��B8R��l�H^ ��0?R��S�j��dgR��+B��2����-,4���F�����ڛc?)Y�I�՟b�0��5�<F)B���xm��bY-/^��H��2��l�
�Ɍ��Y�J�g ����@�H�<.S^��7�1&2Vr��m��ȳ4�%B�m9�Dep�an� B�=[����ɶ|�j͞Ϥθ<< ��u'��	�ī�:�3���0�Y�_�x���MT�]��
_'\ݯϚ,����u��AXN�d��q�+۳���� :%����o��u�~���C%��"?�7�q��*�W�C#XV���^�#Yu�_o)bBqyǮuE6{t9�j�ug\=�4,�=<��pE���|yf9�V��g�(���X  :��=�~`���r:mO�!�v�أe#�	���5�����ǧ}������џ	��-�=οHI��!ZHy���`����M��I��w<���u��ߔ��T���������6�ױ�V9�>F�UT�1a%.w���G-!_����!����,@��>�ׁ�G�OBa=ߙ�1N\�/���ٿ�TBw�o�С,�Њ��c�DGǢ	�@��BQ��P�;ws�vNg�O�'�&��b(qφii����E)Ϥ� ����A�]n�m�v��eY��2m|=��/V�ő�pq�B�Aþ�.���<l��kz�-�h��ȡ+
��spCc��;�j�@Ƒ/'X(쁭�>Dp�q�v85?��%k�ԯy�,��v=G���~�ԩ�o8����F�k�@��Fs�PQ��h���9��UKѼ�O����Q������TF�X���yl'8�2�"e���z���Y��&�<���T	��7(f���w)��=I2[�����Ds2{%��Ƕ��>����cM��{�3P��D��;4�Y�S����&����qQ{���Az<T�ق�=�0�����-�����n"�$�X�:J@|��F3= (�G�u��@D�����+>�?`	(BU�>H��94{�(�������<�,CY$ZbAè�z�����t�0�%�m�@�����ǡm�1���rs����,�;Y��`�Irw�l@B,�^�=�żצ8�G�&7� Z������,Jr �Ũg�rM{!r��pQF��1>��q�`TFZVJ�mr>�-Ki�ն��a���BR�9L�	�P�n�X_J�
�Py��!��+�h�=%R4ǈ�-��Yi{c�
�L�縉 R���Q����(��/�G
乴�Zt�-Gb��$"�>�k�.�8�sφضD��_�KH4>���0M���$��s
�go�9�hm���("s�g�tI�~��¡<8�̫Ϙs��}捗Kg��K/0�@�cj��x[�jv�9�`�R�,9��-剮J�q��LZGZ�����z�- �w���a�p`f8�knQ}V:i�z�6�j�)�C��	!�[�����C�J��Y ֬�@w%���r3ި�;��H���x�������Wo��ʖk~Ww�m"����1> ����UA��14����Z�\z�ڻ}:n@]��@�J�ԈB$� B76�Ì��,�1&�~��Ƴ� Ѯ3�Z�QBH�I�nuܬ�c�!�G�˞e��ن[�N 1j���H,Tʲ�v��*��gV�C5�0�]ڦ~s�z;!�����c�dC��H<)}�*�F(0XD�5��h�^�e줖5�֓���O{LY�Ʋ�O�����R��� @�bυ�>3����l�-��/�;_�I���ǮnFP�xl�v�*�o�8�%��iͭ��z��i7�D��FU������EWd�������������-F(�i�|����0��B=8E v^�f��`�w�O�!/��,K�n! �VK�χ�/�5!�ns��l`3���dm#���m��Ejyp��)W�q@�Zp���������HA�	2@�*A�Y#%���p�P�޿�b�"�O�i+a�]O�t^�2Xr�nS�%S	����j$���(�Jc�
��1#�	��	D�!:v(m���ң�)_9��K������)� �x�U)&�P�
��X��t킁��U������ET�g�t� ��;pM2���Vҟ�%���������'is[�a����e,n2���Z���+�>%����*qIX����B6��cK=�ݹ��4�Ǿo`�:��h��7�l4�����"��I�H�-Ui�|��)iA��u��˼�=^l],�'�Ɂ��+#��ЫB�&[1�S����R�s ���/�&r��R��4�D��.�1���{T�"a��'�Y�=<Gj��t�][|�2�O�p_�?��e�k�u�Wx /�w�@7����p��+�k�,�j�MQl�����%Í�~��v��CY���`��f x����Gm�JX�x˃,��	!$e.x�u1(/ζP	����O2D�.}��23b����JS��;���I[jyB���M�K�{�NV��hSv4��D�W��v��@6�,��z;�VE!?w�Y��\p	�1��e�����ȴ%���c�]{B=7�8X�cEvg؅-��P$�������c?hoK��fR ��_)+��I��xߒ��k"�m�*H��l�{+��^�����;���Y,\M7<���)�*��%���#P:�-Yc�q���*�QG�˲��^�Z'^U�������$}HRt�Ed��1��E�������P4�x��z�̬�f�f����.eėJ����P
�Tq1�dn�VJ� ��&���o���ϼ���SτK�r��:7�0л�y �L�����P� �_@����PR3P[e�W��ٟu�RX��$�h,� ����y�:!*�׹��R���J�	}��~�n�^q3*�j�U fn����R�k��"ŰQ��7�:�y������Zw��;�"k����K&�7q��������flE=:���{�a�����zX$+z4��Z��}f��{]>?0�-�uk�}ș����h�0׹x|H��XF�����#&��|qѴ׋���_K�� HS���Oa���+���8]���e�lԝ�ܚ��
c��Cb�&�}abcT.��^�暩�p'*�v��o-�nFA���x$�� ���"����}�@�6�2�]��������ȩL�l{(�NϮ��G˒��}�?�΃���OT����ӿ��j$ig��w �cn�#�L2aݒБ�?G�mV��,���y����P!���'o�v��i�m��?F����!�<��v������2��f/R�\S$
�G<��RT�&ޛ��*8(?�q�)�kK�"�8Z��
,Un���(��euᏸ���������h\�բ�xI��ʪ~�Fk�YG�w�c�{�>�*�������͖��%7���ˠ��3�̺�m5;v�9N�
`�O[�$��W��,�����mf�zo�����%���:IA��A/ǝ�U	�di���s1����uIпga�p_�`��>�1.	��I<hti9ׅC,���9j��R�F�n��b>�1������[@��p�ren�X	<�l�Z���]^7UV@�~�PC�`%w;����D`�,5�wv��J,�Sb�Q1�,7�r�
��U�����s�5���G�����*��h���|Í�Q?�D�̥0�y�bQ�O�(�Qvomhys��0�!}�%���?#�es��ҷ�����[g���h�PG{d06�!����Gf�Rq�i��� �����]�������P�bO�d�=�����*��@���0���H��]�b��[���s���e�9~��%W֠ ]~����W���y��}�O�p\X��q��x�Z/M|]�&�[uc�Y�V��ǈ�f���E묟w����zi� ��)fx�]Q����=!�E��l4B�@���Z��Iۤ���形1;�ו�U��VO��Z�����i�G�أKm"�g@�1�b���hf����SK63e#n�BNc#���Q���0�k�jU��4����ĤH�
�N�M�F%TTʼv�~����� Ŋ,I<�����|���vGw�p�C ̲�_\����[���l!'��9'�C��\�x�M�?��N��c�Q�[l����aڀ�e�Ǚ��)NyIdn���Yq�U��n�@ ��e�ױ��CH��D�O|ʮ�5F=�z��!�r�}MF�Q�3!v푧����8�320F�Ȗ��-�7حs&|;�3@���(b9�ғ�L3؂���8+'�Ew�߬�g�t�Վ~����7
�cJOR���I��cr�~�KƝ�j#��HhՕs�,�A����������QCO-6�Y��z��$�Y^���=TUj��L��RW�=���_�m_���w��4!i5����kV�-g?n�8?�'yVc=+�d����
��b�K����U,4��AW����� �0���f.�����hx�0ks��%�q�^���w�����r���ر����2���FJ�V"��BSв_��� I+Hu�# ��C'�V#�΃^�B��=t-B���1/�#��{N|��J�#JϤ�r{?(�`0�v�����=[7[fi�������RV���&o���f��s���`w1�@:,��m~�� x�;V+������+r��`)��Wf�Z8��y�#:�Z�%Q[3R�J1Sɳ��{�E��'u�b�
qS�����������T��f#�h���,o"�^n����:c m\����S�]�'6�:2�Dਝ�e3�F4����%�4�zs�p��\C.�y[c82�\�ڰ!r]R���'cp�յ,e�4��N�CL��d��9��y=lwN?[sB�|�~�r�