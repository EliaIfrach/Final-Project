��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��-�ro��i�����/L-�U��lOjj�l]I߫�p3^������_"�'j�ʬn�*W�� �a��;��}���������)t�X�|�r|�~U���;��k��2��%�`�	�c͜��d����/�OB��*$�K�[�>�)v���������~$�sF�]����ZP�6͝*����ĩ�';ɒr����YU�|��#��Yq���65��~�Mduث6z\j���4���E_w3�Cن̷����o�I��Ƃ�G���~T�VO|�θ.YW�9�����I�0�J����r�=fw 	`2K�$]�NF^-F{Ux��L.2OP&~����k2���S�BY�F���iG�H�E��+�%h�<����I�[��G/*/�F��➳��nZ�W����Y�o~r��_�$��\����f�M8D�o�OO���"��D�_U�@��MC�`��.4W��ف�O(��
��,-�h��jn<;���#��'>�鑩�!i����8�1	ZB4J�yY����p>G�����ٯ�`����?C��?��=Y%!��b�IWx+����Q�XjD�I��5��� \�u�u�@n�X�gs"ݚ�i\�X�8�xt���'� �� ��\U,��P>�Q}�������g�]�JJM,��𺪆l�
��z�G�+�QeE"�<���?�PS��"V������FSh�Q��p!�o���M|ln�P2଑��\v����7��e5h����p�C�M"�-�v��4͵ȁF[�=0�$^񗪏E�,ǫ]��e|'�\�D ކ�8{?��WQ��Ж�1ʜ/��(<�n��[�Ú���Zd:d��Oq0AC�Ӭ�({��V*���
�B�n|�ݠ<̕僂�&_����|D��-�G�Y���b~�E�T�J]L~56��� G��������7҄v��k���x������ɨQ�±����8��[��誹�b��ji�XP$����C�GA��-�"�\mEe�Z���	&�bS��<W�N��\j!��z�jgaaS�?������xڟ�:�Le�C���J[�s�<֦i(*��q�(n2f�n�� � ���	+��`���GX?FJ<C5=i4W�v��1�]G}ք��]�A��v��5'��^>k7�V3���"�a�� �B��򁲄5�>s��Α�f��c�wO\[x��B`�.3����U�������X�z�a���i���T�����H{����eUVN�e��$W�R�e�Pө̬�)�"�]6��,}X��Z���vZLF�Re�rl�S�e�7(�$%bzv�$�«d!��e5��6���`�PX���#-H�JjL���ȁ%��\��tI�{���K'�8TQ��,$ٗ�G`�^ë�^]G�Q�_*G�
o�:u��D���,����N)U˧-Ʒr rgC1����0����ɿa
��v�vi�uC ��i���+9B�4���3�����P)W��m���*��ҋ���Tp��ίI�R����\ٕN�[c��V��L�"s�E��^7.�e�78+�J�Bu�XԚ�@�ۣ[wU���V�Ʉ���O	"�,7�����ܯ�����P;?p.h�+2a��mâe�(�W�y0��S���WP�.� U'!2�#��7��0P���p�6F�5!7�&�M��,Sg�b�\w9)5���<�CLa�X`���T�y-��c���E ���)�M t�Oa��jݱvjBb�j��2)�)�w��o��-~�3�H+҃c
�"�>�v��~#�A"�r !tmVT�0�uX��������P��F�	󟶤��v���+d�]D�o�;N�4��}ѥGrZ�����X�	{Н����CⳮK0�i���N��ڭ�?/���~!E��Uu�1�K7	�<D��Z�-\Lf�C*��Ԏ�8vtU ���ă3mv`!695�N,h7]����PDX����_�h]醊�a~�T�����6��pD����~H�PQEM\��7�_��v��U�j��H��\�k�>~�sx9���P�|[4��M�T�h������=�Q臠��?"��*K{�֢�P�fy�����&[v|�۰�Ɂ��LQi�~�%;�g�3l1X4���ʉX��G���-,h�J���c��A.�ܲ�,�@]�ӈ<�ӕR�����%kS��)ঙ�BlJݗ��8�wr�f� ǘb�#�Ҷ$��,�od��W`����cY�
�����rU%��&>��D�p.�]���7�����"/�~˼MRяn<��36Ic#C�čB��'mr4#���1Az|�<��`;��eS\Lh����DS��L��#����$1DW���Z�MHH��
�����3�^(-|�,������WϺ]kU.�|b}?�����3"��I�5�#Suή�Q�!x����nzq^xH%(�l�G�T�%�K(���ZH� y:λ�����oV�إ~{�
�ː�2�L��n{N	�Ē@�:o|�+����y�LP��)*��X�Z��b{����aVP����c/��wK�Ց���O}/l����.WZr��i4���6\��^k�*h���
���5���}�~:��4�;	�)8o��8�ֿ{"(�P��� T]��a�wO@G��G�S3_��b�.��!�0�@�x]Ѭ-�F�e
�Id��{ �Oˋ������sbjX<�ADɖ��닔?�����_��=���hө�7W[o���{��r;�x�(�E�y6Lt��#�T)g��G4����ks��
�%ǂ���>�@Gl���ҢN�`z�N�h^�:A����ae�Q����a7���iv���,Koɬ��۪��o/d9�j]��t�[�{.]�Ԑ�l(��8��us��S�ԴD�s���uM�C�q��G~�9�b��Q�t�	ء���*�_�����Q�,~�.�o�B��6�9���q���"�袖7�6��[%|�|j���}	�NҖ;!E+W�xT�ϴ/��r���@'�	��N����^�1"��x,_�����Fw)-��.إ� "
�_��Im����Ԋ��t��MT=)�����a�\QUQ���2u�o��݂8�ݵ��kC��3:�fA�D��V�ս�����F��P�j\�$�u���`��pD�I��k��_�!�_�ۜ~goy�1�z�Ջ��uȓ�Ce�9�2��%�D��L.¨��
��"�5[;M]p�`�W�#�Q��1o���6�(��3ݶ�`^6Ps����N�[��@�2?`�4j�r�0יă�s�����4���DP��Tc�h~�P�xd#�M Z)1�6���LS��J��9@u�j�
�u�`�I�ˏVT,�b��@�۝��,���Hý�~?�ε�B��ZJ�:v��G�˭�y����y�| >%�,�<<�C�$J�&#��i "�>�@���n�~6�����|R���ѓ w��\=�R�^��dϮ�o1�������纩���f�51�S�-��3�B0=�c����N�3W@��F���˧�	�Ɋ��Y2�1P��D'�Ϫ�[8bRC��2�D J�_�M�lYI �.�l2js0��aN|���ا��T�� $��Mд_c�:*~]j�:�-`��w#��������e:D��(NR�r�;�B�l#��L�����z��'���0�6���cM9[e-���S�z��c���d¾�N���BC�bI�_-H^�vD��ڐ/�E#u���=��)�2�������X79��9;I
g��o[�	6z��%�����и]���t��Dz"\�,�vU'yЁS���U� �PD!qO�ۯ/��՚�?��d�B�s��h�h�n?����r�0GS��30��c�x�l<5�/���}�	0%0l;S�����@���!�J@G-#��'�r��zȿ����,R�Z����.K��C2�:W�a��$e{X�@��Q]�T���"�'
��۽��jت�wR�C�I�;]J�}̘��/_ ���!��؂�5R3�{��A��^hV��%dĎi�������עЪ��6�g�-��b�Le�A�PKB����4�c7�8����=�23DR������VO��x�P�{ܴ;�o9[������y�b��Z�ò�8��|���w����C��Y�����[vj�� B��Q�yr�umk������RM���m\��v�~RH�Rh�)���FF�9���a�zx7׊�����%
�V�|�v��Z�o'������tu�� IX�И�V2�ѽ��Yշ�B;Bcxޟ�e%��9�YKmd��2�P�u�3~�� ����t���w΄r�~� 0 ���%�7G�9$�&���+��b��_���|��{I]��I�j�K�oִN��j��Q�a�j�
 p�)�����dG�:�^�J�^��q,]��Ϋ�֌��Kk�k�J�N��\�8���gn��:0*,�+!n~;#�2i3q�I�޾֨���W	9��%%≾0����n"\F�L�Ŕ���^a��l�(][D����N�%�]{���� �l����(f^�cP"hm�4����^`������՜���^#�hgCp��3�}�2�C;A0l�z� }]ظ
�
��z���W�l �g��v([���Z��a_�R� E�n���i��-��Z�M�Xb��$��U]3=N@�YO� u�#�V�����#��<����`�[�R�sUp2}�?8���&Q3x���Ćn1�G�U���-_�a2��қ|��R���a�H����s^�HE�,���K�ᠷ}l6}����M���ܞ�|
�����6m���EQ���gw��,�Kb���fuz�[���XzRr���)�������s�����Lr]Lr��(��P�h�����T��W�����R�B/|N��̨���v�=�E2��(����\�>M?�vwj9�e!�(n��3Q:̡�q�NŬ�\/���G.��7�A�E�W>�]m(�O��q2�E$?Q����ԒQ �Дq[�������*���_Z:�P\���CQ���1���Р��ks��%�eh�n)	�(E_�驷-��NR'�j���hl�1��cH��C�D/]���&k�������5[y ������!rA�x��g��i"�0�o�����4H=�L"�wt?߾j�W�dNG������f��%�iZ���-�~��f�W
go�`ˡAPQL���VW�x;N���� �e��)��7�g��w�9'���L8�弜����l�Fs�4#�&�$(���n?�+���Ϯ�ʚ���R.K��K���?T6�nԩ����@0��2X�+�>!o���@�,;Q�2{R����ۧτT[�COLE�Ok�����Q�t����X�yw%�[��m�/���0�!y��
��[�RX��sp�ø�z4GV��5��|�(Q�X̠,b2�qC�E����bXcZQ1��-P����v�8��b�+�mс�EM 5A7��T�0����՟[�[�������\$��z���+�t�������iV��y�w�����Hg����sz1}�
�xzd��H��Rt2��v��K��t���X��"�,Q8?�z��TQS���Xο��v?����c�5l��c璬G���S͊'X�����@q��?�m�
�[>� F,�ǄQ�F	E��!�5�>�3�)�5�����Ƣ���z'��������5��ʨJU 3^���B����A��2��s$�����Ԛ93���P�&�y/��� �[|G�g&��z^��Jl�xXw�\l���s�	݆��xW��=��;i�W��s��T��a��$�A�o`������=�Ǳ�wk̐3� ����c���4�w
��<�V�"~�F2�;ޡ�:,CInh���.4 h����gp�P=�|?��kRSNK��QQ�s&$�7�Z��l�]����
�1_�Khу�nƃV�8<zM���]��2�Ot���)�ܼ>����=�0C�V��Ɠ�[���ۛ@U�q�SVtj A5*�Tm�֕8&�m}W PX����1��6�í�U�����$��f&x���zPi�?��5k�ß���/&r0M�&Y?���93A�w��m����Iܬ��\3k�{cN��������!Q�ټ���
��K��� �	�;G#�������Q���׼*x�j�zZHdkwO;�r����~-���>�=��+��?�M��7�x8�����V��Z�{yEάA�\���vA�~!fY�?��57�85��RQ��a�mW;Ӥ(W�#���(�B�ӗ [���&ή#�"E�(�K@��0�{b�S7My�R��Ȇ��XQ�(3aIW6t+6�3�3��<� ?sV)*n�]C�GID�%�qS�K�w&ѯ#S��m�>��2��c�3�\S�h�	� ��Q��V���o�9���ʒw��"/��b�a������t�y���^)�<��z�����9T0��hC�p���u�4�b�`����6�v �w41]Tк
�zA�bp5�L0]�苁�����\lPdq3����[����(���|��)������a.#�a��'�tFSr>���!5`�����W\�~�����m��W�����+�đL��E&���W�	������G�K7D!q7��+"� �BRSYX�z�����\	����t=рo���~c�#�M~��e�R#Pϯ�5$7:Z!��C���G '���)��E�<:����3D����b3"`�����WQ�)���e�I�t%�&���B*������o7�m����~E(*O+6�EӃ��e���!k.9ZF
DR�/��tU$���Ʉnc�c��(Q�+6����z�l��g��>�A�OIo�!Y��s�Qd�Ȉ��-�NJ�=7Dǹ��i��B�D��,�]�p� Aǟ�ڮ���� Ӄr^�G`��O��a�=*w>�2j�2����W��Q�kA9|�Lΐ�#O0���H���C/c��e�y�
 ��8��>Ό��+���`:�+�R�1CrB�CF���8���4����Җt.t� ���I���I���X�/uщ����gV-W𶩖4ib��������F�!�/�酗O�b��Y�֎�2��kl�J��$�G��}B��l*�t��7D�+0Qd�a�~ ��j2�I��_��D�A��ְ��"C?��䪆�{��e�O��bH����6��):�ix�y
CA�w�o�8Z���A���ߺ��3A���a��t������G�����y'	��>�*�������O���9��>d�].��6/P��C���!�
�B�l� �i��N>� fU���X�6������fϊ)$�;4v(o�,T�ܾ(%��� ,OP�2|]s>B�Y\w#��)�"�����c<�Aa��}4�������}&��E�C��S�������h����Φ^�)����� �b�ׅKt���":�x��l�� MGd�<
��ЦG���L������HZ|oW�$i$����PؗO`;(��u�6	�@s{A�:���|��$Ub��4G��&#|B	� ��p e|�O�V(T�0�1?�� *U��^�����,H�7AjS���)Yj &�B�4�^B���V����5��e�v��#�P�(<���]��#ow��-Ə ��Aw����5;���K�}ﲩ��:.�rf�㴯���u��_.�����dk�e�u�HO
W{>ið���<�6A���� ������������K������L��G�2��I�ȉ�1-vo��:�L[�����=?�.szqH�V�SD\��;E�rǚ�)6�U���|��m���HL���˶��e�l�l����.}��X�a��S_��ȕ�U�E.7�_^��f�Ȫ��ё8��?k�i�@9t�����þq�	'������!(�{��Q-�����>��i %���|3-�	�!�����V��C=*�zb#�4����M-������#�*~h^��T��#��{{n|���2����� 2���S���5���f�Ve ,AH�*�Wĵ�B��	̦�\NKy���߮���%�N>so�������1�>�2�&�	.T�F�޲��9P������2E�i�����R��ܢ��5�9�
�)S����7��k�$���_eD��%��6��z.мuLU�Ǿ9rFf�S�G�l0�ʓ�Z�
���U_E�:K����_j��!7�M�TxX�	��l�����0�)-�^���9��._P֘cN�#����*A��F�������vAcT����x}r�%ߞ�:�ܔ���cQ�H2O^o�I��t ��[ћ���:��2��ۏ�%?Vȣ2K�x!Q�$���5)U#�;�Ֆ1{Ex���0��8?��^Z�Ԛ���o�U�ؘ��<��O)`ϲС����(&.qC��&t�:��z�U�x���mA�A��P(��* %,q�Tˊ�g>�3I��k�\ǉ� ��K����j*3L�6Ͽ%'{�s������Y�%~����:�ɐ�7/	�%c�E���9�#,ĭ������'!�7E&M�`b&ҩ�G����q	�<��j��0�~.�D�.k�0ZfdX}I��k��E��@�˩�=��+�h���m�*.�#ثb�yS�u��?�zA�Y��
���>�@� `e�:���XH���/�D������(z��{�=:�^��XH}�L}�{p+��4���R���߃N*�ŀU%f��;�/��ķQ���k1�g�ܴi�Y�������Nf�߫�u�V�b��<ۺS��^�;�Ax�$;���J�����m-�'Ǡ}Y������T#o?x��`�l�$���N�F�>e�����}¦��
w�Y,���Q���	,�#-�q7�L����7�����'��;��X|ei�����aGS�e��-k�������
����Z�݀�a\
���&Y�T�N4����H�j��N�߼^��z7�G�bPL�����5Z�]����&��L2+�f3�wmu�S9L�bc⵴t�d ��a�z5fL`O��˜/
�[���E�%�r�`