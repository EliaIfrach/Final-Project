��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
O���w3�2��P�?��}�Q���)�;��L E���,�ڬ��ϭ�w>�A�'āb|�}��!�P���I8F `i�q��6�d�V0g�B�?��5�!�WDc9��"�\ӂeĊ|�#'�M��=��,ɀ"�0wCQ�f)��>��q��K�'^bq�5�w�dF���&񏥲�Ǐ���{���?
��ؤ�	��M����Yu��~�</�d X/�%�
J~Ql%��9"�ta�e5O�%|'�����(����n���� �E�:��.o�Aa8��V���f-�C@ q�j�9�<v���ۓF�Y����%=��8Kr��?:��� ��m��0�#}݌H�C�zǑZ�K�Q[y��d߈��?�H:B�uU�w�n4`��!!��B6f�t�����'`?��gv²D�l����@�e�ة#�ne�8S�[b�BeaM�+T:'��Ϭ���b�L2�Z5R�����GLN��[���)4��J����U|�ցcr�����^7����A-;�˳/uԉ�PU՜>0,7�\�]D�����ڐZ�B�&��.���S{4�Ǒ�c��/�B��?yRO	�{1$��J�k�A��t�ⵃ��T���K��o��V�bc�m���V+�JW����nW��l)�մ�ih�3����,ʈd�a��˘<��@n��@V�<E_��;��{�}>jo|(����ފ���o�"d�U�����L�{�w�YIxM1=��1,Q�W�kH�]�A��q�����\��y����Lr�`P����ue�H�O~�sU9�X�^�V ~e!���@[��vmUR�E��9W7?�4�6O ����e���K�VK'���7�I�fc/%��5�Á"�������J�@���2 R#3o0+��6�Em�;�=�b0F�z�7�h"�΅n׹����I�
"O<����Q8Q^p�(AP�uCSj �f�p�/�nN;S����G��1�Lv���1jm�3	��ܵ����`�fB.T��Xo�׏����j��W�^��`�F��l���GP}|�rEQ�H��.3A�Z��k�|!�A���DAy ����m鷨�]�հK@��#)�c��]16w )�712&��8�N7�B]^=�%�J]����@���S���Quwwv 	21��O�r}��r���-�cS��)���:q �tx���F�R����H<��&4ζ/&.~3�֨��e��;�fb7�&���m/�!�؍�<EN��e�=���j����n�K�Q��W�9��{_�XF���P�4��Q-���T���t�#�����&��j�B��r�H@���*��.��]�{L�E�K��!\z���?��5D���+�L�
=)��f����^*�N/ٌ�c�����������@2�G�o|�{���	������(ޮٴB�+=��i�@
6C��h?[�t�2ݬ��%���k�1���l��sh#r �����/�Wu��훀��J1d=��K�5�Ȉ�'��5R9�$l����;H�ӮM��e�/>���ˏ�X�E�rbd��t�,�[�����>��7d��/�����D��3������:e�D�ݜ�?c.;u��M_��c��+�Ưǒ���	����v-��H�w���o��ۇ~�yh�z,;�~p���W�)��*:�v��O�|LL[�<�j-Q쟧��?Qd����G�;Tծ�����t�e�A�f�&�a5��������j�D!D�'�#�>&3~�y�L�������\-ݦV:N�S���0���t �H\�P>N-q���*2j���w7
�	� !e&#!��.�d�S�ĻL�|t�s{��÷)����M�?�\F��*����VC���l-�_dB�D�</+�moq�X)��>�H)^q�p&��y�ް��"Q�8!�@<���E���hU�@��~g��ʥH�V^e�t3W�݆y�\�?s41�m�E*2����� ����<�|������'	��(��:;��=��b�s!r�7��`��x�*?�Ep�e�@aEuvD��y��� Ruv�Q��As%q�����D��u=����P��@��Gnc2���B�p�V�t' �Y��7����*ڈ��G���6b�g����W��8���3���W$����l�H<�m�d�7`Rtu��;Y���}�)pH'�A��&��+�Ѹ.;�
i���� ���<���:#������ʅcҫd�a�s!�����t�f�M��\Fi�~�3����j���Ď�6(IOVe��=H�wѾ�*���l�#9����d�T'*[.*�S}ߞs�q����&˙�^�+& c������Fz�{�!Y��Ț_0�1�j/]וƴ���cj���e]&�@�=4�Y[���%G���Ig	��7��;t�v�c�ƕ�w�F�?���I�+�X�:\����]�)	�^YO�n�{F�O��nSD�Gv�}j�o3݄�5��ׁP �&��bY�<e;W+@�����~YT��I9v�w&ȑ<榾�i
U�x�*xÓ��6/.�r����K�0
o7��/֬����$���,S�ޥ\�J���T��Z����&;�΀�����!�0z^�d%v��E�������@Jk�l���������nU織����"2{du�ʰ���;��d4NBJÓ��jޘ{�8�v''�؅RZy4�H,S��4m&���z]���&��3
y��ح��K�YRx�'�1���&���O�*�1�L���<C�A'ϧ��3�I���B������B�~Hyn�n��o��ؕ�BpR��J���&�3�>�2���.���5@6�/�EO�ߊ�T
�"��|�=�אX����w4r~"G�K�<�v�7p �^�6E~vmԼg+�J�A��r���l$;~��T�]֞
��_�̘���f�~H�S)2~�^7�Okl�v�׆�û�44)*j/���(��u��Q~�쮮4��L����2{�� f���y�
�����G�����\�U�{��j������Jؗ��Z}���:�[M ���G��>�K~�_��n�0c:�� �|��9���:�YMB�O, ���I�6'���j��p������s���|�	�*и�NE �o[�?�yu���@��e��[��B8_ �5V	��ڣ�����	�/u~N
;/�ktAu���%�t�/9��G?�PqR�o�j!�{,Ѿ����ڱ�!����2���"P=˕�Q���Ȥ�ѿ�P�!yr#�i�����T��/�<��2rn>ٳ��1W>H�g Ow����g<B�:_4�	������A�