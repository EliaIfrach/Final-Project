��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A�m0wS�֧�e���u�`�4�~�8_�E��r-	o�Bћ�`U���������ob5=Z����|�s�-:�r��';��N�L����;��½�P�.3��y��/���lU`ӽP��ۣ�#+��og7I���ʞ�V֒/tB��X����,�@ҫh��@�ZX�
��ψ��S���z�u5	�9�h4��g�q4V%Cz�9k�����@�_�To� n��(���ʬx l���?�2�/����Ȉk�H{�L�C~��iT�|�$<k�;I%g����0�)�.fB�dq���i���FN=���G���$����uB��+D#��2�����:Ư�rn""��� C0O�N�P�'��i6a�7����dG��S�Y��+A�Sg���Aׇ���[�~�_���oII��u�/K|�i�oh߽ 9]���h�@��R�*� g��lc��s�鶉C<����L��Td�d�B�����K�[#���Ԟ��d��sO���9s���a;c��`qKͻС�#9�o�q�g��y��?E��\r݅�m�����<I���/����;�o�x�{:e圯Oy7�H
�9S2��k��*V�+����3���5W�8$���k��6�{6X��<@�gz+��; C�
x�f##3��n�ו��������q?��wb�K��2�yM��'+!���R*G:y�"�YK�n��w�O��r#�仸܈��{!nS@�K��T�+vPaeL'������XG�U�]Fm�U�7;'�'Rs�*����/�}�ոx��K�"5��7-�����74q�<�A�Q�Ffz{�(�*��Վ�.�.,�����U*r~�8dZ#u/�G�y�T�dXBr��ǉj"��G�8Y%���k(�+*�]\Q/ׄ5�����^�+Ś�"b`ӳa[�p��.M�~n��jt�����Iް;���p&��m��d��m���+�/i�k����V��.T� �I��m@��M:��|�~�����4�6�N��t]h:�˥�S��8���.��l�($�n�����
��f��?���R������Y�[��%�����T#@E��XvzקV��>ș�&�¸F���\�F��$�����b�E�]o�͹�⏪�m�$�����[��U�`¡����L�%C�!N���q&SO����8�\��ј�0S6���9b��9|m���,������Ȩ�T�0���w��jN9��%�s$�l<���~'�$�;ά]���=yN� .�9D߰:w'oƇ��`~]zm�������a �U�M���?�uƘ�L�c�6m9�b��bä5�����R>�:��H���4FW���癪�Kyi����G�ttf��P]�l<�K��}1�:���5k�s�-�-rfnP��(�-{��_��q;%be&�07�c͛��𒚍3�~��)D}��p_����ZQ�{I\���*���6&�SH���#��+p���&Y7��C�=7�'�rj�@���}s������`��i���O^8�G���ԫ�َ]m>f��j�vƮZ������!ʇq*��Fp�1��~�NUtzuۧDz���eY[P��"�xAW죲O|!�n!�P��f d��Iܓ󏥇�>{�r}��B ���^���u�<Ilk�7-%�G�O:�k��/��t��\_�~��8��^�y*���cc�Z�Yu+���N�x�254K��惎tW��T�~�밎��(w��x&Ѻ�<ظ�V�(��GåMC @���~���	��q"S"I��������l�z%�@�.�H�-�����x؁��UK�I�i�0[pl8"t�7f �����H���σvsm�t��GӶ��[�����;=|��h���0;z~96�{-����.�M�>K:��jե�%��xE�g�������h����h��J�ZϺ�"=� ���	���}���,������6��L�ʫ�.+Z�(Ie�9ڣT��9�o�G��tF�F���v�qj�½�kY�o���X��f�nӋ�4�������NڤZ�^�?zm{/�lA��#{���8��l�{.��>'�zb9h���Si�����Xi;�tt�,�E"�4� f��pm�xD�+����~1v�lt	�vnҶ���)*���(,{�x?��]O�@�%{�����v���2{�?�4c�����Q�EMq��5�gQ�n!�ײ�1�H��ԥ�φ5"�������Q�q~�}��"��9$KB*Hî�andQ �Պ�n�+��+���.�B{giaO�,`�����?��vԂ���3�Cw�����]����,�ځ�uq��m���@�p����]\s���'C�}�-o@�o1��]
F� $� ؑΔ�����-�؈y���$D�w9�"V��#t�]Ұw31r�;G�W@[u���:�9�j���<B8�_?��<��Y����SWҪT	UGy��tל�t3 {C��=�66��[�"!��Y�w���	,�I�3g?,�\6�ƻЬKƎd9�(�߳���Qr1,�R0����h?V�+ŷ8b��ҷ�D�?�~��5����,�NM:����	�'�' �/�$	�.����"6�e�;�h�w��LX����LRg��杉���������d��;"-��ӓ\dBd��@Ot�]0e�4�R.o���'��Ɛ�ҟ���t�T��X�Su}��H���O��.��'�s��l�h��=c��f	\��H1u�wY�XQ�T`Zs1ҹ��w53SO0pyX��J��Ƣ�+�"o�e/H���ݼ�o���%ʑP	l����㡛�m���r���XD�\b#'RD��DH*=�|� 
]z�%Z��� =�:,��Z��D^��mS����U�GEe�/��U)�A�O"�v�ץA�SҴ�T�����Td��e��W`36����yFʭ��&���>N����`�NT#��!���R�%˰5r�M�B�����.�XW:)�4��	���_�e�E<�ra�&v��{}�EԦrU�!����y�|��
���I��2���	�:9�Sn�����CЃ��p�k�����u�x~y�{v��>�k�Gd�i�_���<bRS/ &�D��:�k��,�_MR9>�A��]]�3��%��{oAH^�
�P!��(�s�u��,�-n1k=��i~�.�����z�s�����Kw�!�s�>Ӽ�$�CU���5�9dE&(/��^��F�j���B��!�p�>'���T}4�w���I�0yn��l�@�'{�c��8u��(�X�-"�"�c�?�'�sɋM����>�$a�M~9Gj��>ں���[��t�[��!%���.y�L���{ޮG���iln �UK����y�e@���q:�o���)��)���{�(�|���U�ܖ��c�^�p�@�T-����i���M�򒟬s�q�M��U�_L�S�ø,��=����S-�!�F�S.��=i�i�L��z�(��x��Gj�.Iy�O�.��aP#�| ��{r${��m֣R�`g��Q�F�7�)�si�������!/��.w����,�;*�-�ch�Uk5�k[S2F��r.\���ǯ"*��-���3u��i��?2��V=��3��T8��D�I�9+�I,W
��q�]���ǲ��˜�q�x����5xU���ɒ*J��s��dk^��&3���pչ���#�,�a�˪+vs�RdS�XD��ı�z����杘ھ�&�h!ԳfY�Z�d���Cd�О�h�i�Jt��b!v�F�^NZ��X�?�R�r���n���ed {�f�ۥ9���q������_��	Yn�@��1nY�F�;��������������y���FrS�;�FU��āt��S����j�v�6�?��g$G[P]���=n�z�_s��Y��.VQ��m�r��C�zئ��ރx�A.ղ<#Z���J!�� ���N�y�e� �Of��6�7 ���U��ɶ����[��}��Q��e,o��0�����Aη+��q�۠��k}��HE���42'?�	�����%���WJ?�K]͎p�c����! Z���})�e�"z"�aw�;l��K��Gq�}�k3�OsM2��wD�JsBv��T�������ڮ�om��{1�����dN�F��=�K=�;�O;�s�F�T��]�R3�ey5��M]��k���	��~3PR�֙ʱk@�9�;sh�@
�p��#<G�ɿ�z"ߕz>D���|��ˊ�����v���[��h˻m`��;4��#��-�<1�zจ�O(�1X-��}.�y+*؊�jg�܌)�#��7�޶G�DB������0�n��,b��*�2���,erǈ��G m��jb��(�[EФmIL!k<	��oؔ���^��x^�{I�Zu�2�&�è��\�� �� ~L|ͣ��f; ϊ->���CF<�E���k��"���9Ŷ^~~'=�pd{��Ó]�h��$��l�ǣ��Cf��c�pvaJoGv��%�[��ANW���S���dk�/��f(ͅ����-�K�r\
��@� /���l����Z/Y4�߱/�|j�֡����]������
�=zn�XtˤRD+���M���2����_��q��z��ăLC��Pf�5���Kxj���d7�LV�?��$ʈ 5m�����6�; 	6L��h��᫙��A�������O`0G4����0�K�uCT��S���*o�E����W85�L��U}p���:�@��]c�r�J�L�7@
��I��:ނNU�YB�0�q`WD��q��Z|�~a|b{Q]H6�)?:U�w/yH-����E&:�v���1T��:��l�Az�S̬�<2�U�E�����R�Ѥ��IDe3Y�CL�]�Ig�.���K0R������,т3A?���YƩ�I�.�ߐ�x��I�@	���A�+m	�2����i��k��N��ԙ?�Dw�{�R
U?�)���R�_[W���4�H%9����ס"�P��=���M�J��@��ɔ�[��ã�W��O�[�i�8�
�H��X �������٢�۲�?]:|�g_yaf$������\[�B>��/H�_�2�Ǝά5�+@���ѽ���CSnw��ju����O@␫�<�t�B��^K#yDբ�@yr�5���EV���v����\iZ�|9����wn�8f�%��܍y=�MK��r-}�3cOh>QQ�/L���L�=��4FHm�|OXDSmb�,%;k���D��2�0N8��d����74�gOf�ԥ?�p=ԱH��B+6��m��CҺ�fȕ�Nh�G�sl;g{r��`Jb~ 4m�z��tl)�%?rv�Age%Fl�
��EJ�<�3c�bU�%+0b��b�&+Z"PH&��/ �a�UJ���|�}���o�UeϺ�`b��y����̕0�����_܊��6�F��S8�=�J�āN��y<���c|���� ���whk�gZe^�h 2(Z�ڱ�]�:�����c�A�U�<�3v�(cv�#Z���\UD�ڹ�Z&Bu���o�@���``�� Ew��r�"�2���A�����DU����Il�s��
�Jb�6 �`om4�nPdT��O���x%�Q��e��|����ϯB����]$c����u�.e�LO�Ue���K�v����e����	��+)U��b����!L8���c��))!Exx���_�M���ø��$��B���	��X��H����m�"�1�C�W0 h(Ye]7yBӭ�I�
?5(cҿ/.�@x�"dB���6����W���;�e"�2P�\�g��b8�m�1��b@�Yk��Ø���������B��gX�Pan�~`ŜWfèO��aDh/�wr� ��e�xo��|�-�b3_7]
�-p�"�	����d�y��P��_ْ�	��aG�N&QJ��<xZ�e� D���D?�à����;����������V�۔"ݹ^h�����#��&#���-p�^����>�9ͩ8��t�i�"���E=�
�S�i��0TFְV- ��y���c�{�FZ�?�_���^��&�{�/������Ev1�_�i�0����)*)寇REy
q|�1���&���3��%������+��AjSQ����}��X���L.��m���j�&�N7b�,Pv�-�n8�>y�?�-����l�L�����}��E�7���s���	R���P���?��^ϡ��W2��=��br���N�"@�˼ht��:#���GNm����h�(0�%U�FF��m�:�[#/����\	��ľ8���Z��ሠ?�g �R�c�!��v���['L��D泙}N�/q��H�9K���^t���Wƞg[
w �6�6Ҹ��.�[>�n�}�q�3~���v������1*a$�>"	<������X���<�[�G92m��n7x�^�%T,�S�e��*�b�]�x �`Ѧ��=��Du������ZW�ki��-KO�Q��64Tf��������A�R4�����)�n�|���D�7Bm��/w���W�Q��M�Uy����l��1��{$@�ؐ�~*G�Fe� �%D�p�F�⺩�X���A�.ޣ�FȎ�{c�7=Ǘ<�4��&ǁ��W�$L&k,B���Y�g�IY���?j�D��yFMo�������F�k��2��Z�<$�Y ����T�H�ES�Լ�p�1�o�(=�l
;��:��ۍ�z��8���z��w�7�\,�Ͽ�쀤\�;_�C?�K0 R5�׌��R�#�5#�J����zUg��1�X�rv��������}��UĿ�l@�؍���	���k��EuBI�a�c�(+��BA�ڋē�"����:�o�����^�~��3_d_�����I��6�J����#�K�R{��J���#������f�eUp����C-�Fss��J���b�1��������[�	&��Y�)����"ia���G2SB�r���e������_^�Ƃ��*l��L9�$���BN+ ��TJ��GZ}�ˡ"FYV�Գ��hD�+��SǇAI���\��;���Mktx"����쉄��$;泍�Gɯ)$�_(��U���&Z1���U�"v?hc����u�)�l{��|Њ�5�ڂaTڦd����6��^0�7�s߀�FI�O���"aW��
%e+���ILa�e[���@�Aݝ����r2��4�4���G7�����&��d	�%���E�ǔRme�1���l:�H�W6�3�B͎>%e��Z��Ik�v�y)~����50K�NMW�ƴ2Y�����%���܌qb7����Z�(|�-^�y����h��e`����X�@&��Tj:� �B\��^����Gϭ��uO�*�,� s�����U9*�x�\��F�"����I����$DK!��o�6\��V����}+���P1��܀ңeG��
�f
ʎ3u����̹�@e?nm!��1�-��59;;~�z�b*4���&��,�
e���o�j+�'T)�.�*��Ԏa���fcU�*q�S��t�;Q�4��	�s ����7�%���Z�������F�M,�V�d �"op�'�� �C��a%7d9=|8�X�����$�TI�f���}nR�knG��+��v�6BX��k$e��3	��w�6k�!�7N��L��4<���c��)z?`�� n���,(^,#����HY����jA֋�����S��zd��{H���O���h�3�`־N�+��Hq�#m�~sT��,A1{f���I��-�]~{\3��9?�����Z�Ó�S���Q�c&~��g=�a��.����]�!�v���ܝ訷�ޢv �Be���9�k�׹���#PR�@.���\�a0�e�m7��c�������:���k.�P�s�·��ǋ�O���ӛL�wt�ű��Hԃ�;J�U�����O���|�([�TY~��S�����K�_�KO�p��9�c{����}���X�$y���*Ic��\�j�N�3�� ��/����viۤ��G�mv��o���{J����d�"��G\0����؋}��?���^��H���U⃾/4����Z8����@�K�M(�6i���p�{n��W��9Z��J�1��ƃ�0�Z�4���.�۶�s�oЛl�*��C>XG �	f��	 Ϣy�Ѽn�N���j��B�;@e@֓�6�=ϻ?���wD�G�\� ���|U�Xg�soh�y��v�G�6����L@b�:��ZR|���3�o}f����p0�
 �y�Y��̡6�%��'��9͞w�VmM;�x�%HnN*:��^>\~�fn#���4e��1�-MU{�58)�Gs�-��jP4,ۡ1-�M�
�L�q�z���)���:���,r��f�;AJ�q�����K�j�6�j��oqi���?��N��ĸe�5͆�O#.?e�Y���<�q��p�d������<�I� 4��Я�?�#�j'����~}t@TU@Ia|�HW�h�T��^�R�|�^�f�ffJ߇o�7�?_uo�Q8#sOkݓ���c���$#U9(�xJ�i�&e.&Y�m�{g�]s�C��0�7��_�}u?�p+�}���`�&���q�P�ㄽ����x�l���{ˊ�����[s�v��,�K��P�U'RBʸ��,����*}w��!�7��s�2*V�<���NF�YY/�5��J�u�7��,�d(�(���}�,���
M)b@�U�j˩��0f��ſav���b������a�b��}�%<�hb�3hIr ��c-h�����k����2��{���l�Iu��\�I5, ��w�c���D��	7�^U�<�5�T�)"J�X�ɲ��Th���`�E��I�zBG��IW�5Ϲ+Q3��.��=e�ը1�rT <p6�J��Y�5��j�h�|r���j2��v��S���_�ͫ�7W���-\E�W��z��*�Rx������E�/փP�#��E��(�*4�v�,H��DT@TK|��s3�Tj��M�������gv����/(S]�U�:�Vz|ث1�y��eN�����ڤ���ǯ��oo�֧��ܻ�ʔ��q��-�C���0]�� ̌{�m�X%�!x�v��ΐln�^�y���w�� �M2bСf�,�7�������O6"��Ǌ�Tr�޳�HW(��E�z��u�T�,w
��{���r��>����0`��p6�o�s�)���`������r�/��'.�?�_�+c3�L� Q���Z�$]6I���:���}���hl������9+`Tβ�]x�t�+�=���AH�!�8b�<�,����·h:�����8be���G�W�:���*;��C�,s03PZ		!�خ��0�@�]��S��&J��R����Zq*�ZL9�D,)���4�d6R<�T�'�Z�����q]6��84��c��>�D�;�C�9�2�$�K&��u�а5��b}����l�ر��'hO� ��^��b�7��O������~�Ct[Xu��n��8]J�Eo�o��U�G�o3)6�K.K^9@X�l��A���ߎ�PofO	u�� CS�F�|�J�(��6S�)|`�sև�~۠:�P2�/�)�v�q�wbhj�Q�7�:H:�)���)ob��GR%4�AT��zgv�R��Hi{x�y�F �!�� �>�+b
��:����o�k�E6o�,m �F�*b^�i^�5��f"r��ub�6�E��_}���/ԍJ
۰�u�*�X