��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
<�\-���C��ʴ�]O��6e�v�ֈ�}Agǥ��!X8���h�Hۃ^�,S�J��r��/;�!�f��=������������Bp}�����ߛ^�rMM���kb;�!o�������/�'�������}�F�>O����3C�smF���c��}��Պh�p����V2[��~&�)s��?GU����Зa��5;]��`�ܟ���ma�;�<Xv.��p������[��3O�~ދJ�����۟����i%H�ʽFi�S3ѥN�,�֒�&�C^�WHWX�һ�\���`�!�w��惕�#'n�{�S���6����fR0)G���Qw�����3G��=�f�Lj�='l<t��P��V��>O����$��E��uBܕ51��7�� Xُ"��MWYK���ՠ�M�*������ҏ�nɴ��0C�&�t�׿=OCaKV�H\oBږl����+]yF\��)u�V,:�L�x!���L,Gy))g�x\O�Ys�J0�ozx��p=n36��mI����F�G^��)dK���5�z(��s>ɼC��5�y��W~�Z����Pˬ��-/�G��$�gŮ��TE/�hL�`���|,D��`ُy���J�����@��ke1[�q���)z+
h_3=
h��7f�l��BL��N�n�Bފa�����x�]�j0(q��}Xr�7Ɗ�������Bc��d�L��?a�Ѹ�"�E^��4ޯ0�ָD��$9~y�*���BH���_!��6�w�G�@/?�=@���\�hY,X˸J?(��1��M���u1b��ɶ��1"��U�NY�����*撝�Ah�V���}�.�$�f8�*�3�t��s�\^�E9B�b�+[�W��L��?�g x�s\�י�Y��`�����TrQx/���5�"7�+�%5(DF>i���7��
���`��8|i*2�����e�j�/D�����>�yh����K�n��f�g�#󯑻��&�VJ�Ix��Ӷ):O7��	�L��$��[�Gm�rT!�Pa8��
"~���l^�@�\D�fu8�A{
�%/���f=�)n�%dҤ��UU8�g�_ SӲkX�O��#��r��"aF�9��3k�(�p�"Yn�;f�e�0��A ��ϳ}G�nF����W`�A��]���VLA>�y����0<��([�,���S�q�.)H���"6��>-��6�7�����w��%�#�v�*
���ci��<�T��!�#�tܛi�&���J3B<*)��x�.i�ަ���jzM�h5���*��ʫ�
e�O(��F�A�L�h���� ���Dq�hzEA�G�>b��5�j�
O�5�K��I#�.tau����a�'&��(��Q�m�FJVe$B��G�ȉ�8���q�%���I��F_���FL�͗"�!�:�2�W���q��Gսy�7��/���-�����[I4��Ŗ��@��q��3��Lw�����mwq"+b5_���Ty/\�?���=@�U%�{"؎-�c���L�_��)"4���6�Ҷݺ��0�_DE0  ��\����T�����$����( �5��j�`�%��p���:���/b�ǟ�<�����&���3�j_N�g?�ҽ�GȄ[&N�o�Z
����2Ո�( 'Z�ʵ��:��a��˜�t����"$(�}���B����D�j��F�~[��E�����%wyB؎;آ�p�M��Q(���i/�q������r�|_}��Bmo\�~�#{�IE@n�Y�6�c���u5���g�����Ѹ�Z5ͽ����g�t"=����ױLx >�m���\BD-І]\2D��d^�>���e�n+�Lpa+å��C7�:r}z@�2�p���G��7o,�Rwá��6_�7H�GWD�3��O�c�������$'e�v�+iI_b�<K�b!�5��TF�_WNi'�.bݖ�Q�br�%�J��Cűt쩅�p��� +qC��[�ZQ/�����p/�)^͋.e7d���\�B�����1�3-�I�,�m�2x�Hh�/�dG6�������ʅ���w��Mnus�6R�o*��:�ey��vc;�2K=n�62G���w-m[��E2����2��Z��!� 7�����B�W��̫R��!���h��TG/�����,��P쉪1���W<1)^�V �Y��rIr�ά'_j�׃`��"��͕�� l���" �2��r;ҕ�ݴ]h�[9�.9Yt�<�s��iTlcq=��]����v�W�b�rjq���v�7Wk�<��J��˖���`T�;�����b�֡?�����衜������M����N�Q��*w��� $)m��
BF��"؈c�Z���o�=��]�>JF���P��@�J���K�hp�1������2RK�tw��z��bP�bL�4,"�9�k�5Д��s�t|��y��s��iE�禛ĠnH5P��~����L�����d�i���cUB#H��	�j�F�h)-�E-���x�����E5~�LqV�ʯ��!�Hq�v��Ĺ@:o@���]��2�k�RzP	P'���Vz���]��d�R+͔+��E`B_b>H(m5S+�,'�4��K��������U+�LQ�����ƟʕXЏ,�P����jڈp�Ps=���}|���Ήg���am;S-r�L+]�%c^�kR9>���J���Z�yh���3 �mD�������[��Tot�3֥��k������n��@iO,Ժ+L%|���'�W�܀��ցe�'H�l	����r�9�3]����}S'�8�V�|O��Z�KрN���t!�+@r��1a����wo�c3�-��@�;?�����:�Y�����\ ���`'i���ʲ[�5DRꦿ؄�ˬho<l���NR|�p�n2���n��t��=!�B��K�e�|m��s��>�բ3_;�L[�&�PjB����Q{��H�E�'���Xe��ʐ�"m֤ '��\1��Sq1�i?B���]�4\\ܥI_�*��_l��� �A ��z�����?�<2E�)*���8H�
e, �^���i�P��[pM����6ANd�=�Ռ 9�֣%ߏ�U���B�����c��H��[x��ȼ8v��}�<�	����Z֬P$����Void�A�b2t���¼��	w�)w�hWc�ۄ��[�w�Z����bL2���ڀ��j��zZ=d���Ot�c~�Oox� {*�]S�߉/6wE���a@>�2�,�0����0*������ߓ%��s��.��2	��9�������{$��U	!mbn PoZ9t6�FA����uL��x8P O�\B�:k�bh]�&J�캷�!o�;�>��'X������l�@ qdC��uQ�5�������(��s�l5`�w]ҕ- 90zi�t��"��f�y)j�q�VD�k�Q�P1
ߡ�f�5H�W�ޛZ�� ��p[
C}����ݑ�5<d�K%�����Q��\a���j�T�`@�5����\�0:��g|Ӌ ���(�3p��RmN��J�ݏ����ĥi�Z`����	��D
a����/���N���2�rZ���V�B��%P˷S�8�xfցKF�
ଘeWζ�WcN/���4�R� ��Mo��{;��sK��F�gJ_߁��f/��k��j��2$�o��6U�}�e�_ӆ���'O ����0�Ѧ_��~&���uk'������o]�f]3��-��L<!Q:M[e�K|��F��Ϗ����uN P@�����k�Ik�F�.�މS7���� #��{�w{\�91#�h�ë:n��^�KW[�7��܋�V0]贻ʌ<��x��U�4k�f/!}��S�Řty�P�-�[%���
��\9vR3�9�z4��^&`Z��B�v���/җ_�����x|Ή�Ζ����~ ǀ��ֽ��4{S@̘����>��wt=Yz9"/X�-N]n���C��Rn��
��J�0��02u����~�?m�����EE�R;&�X��c����]/�]�o��D_4X �z��ޥTƑ��#fɉ�i��5�1 cџ�P�)�̶�X?�`-.���v�(����1D&�0I�\r%q����ț�gv	�/p�A�WO��)a���~��p�Yڂ��#��
%��	�j���G��NE)�%�[ٮΐ��������HY�Z�I23f��#v}.VN��q����ҵX����a�@�k:������8P�i�n��ӫz~���u�߭�J�QJ�����X����6�P�qʎvvk�T�[��F1-x��S�~�Bi��NLpr�V�	�L��
Y���:(åH�ͯҗ��J���{i��xź.��-fLyo���Xm����5/���An�[�������a�NNUm}����f� �#5�FL�uv��A��G)f�9��JEQH�)�{S{ӑ�z�M�vv�C�X�X�A�G����P�b�b(�~خ���$���ә�^��f��FbS`�x�X�3�-�R�#�f��r eAMm9rPn�\O�1�2����Tn���F,�U�����V'��T�y�[:l��� ��歉���k{�( �pX�"Ȣ �K�؀���b7�"0R��Sr�l�T�,쳖�Y��C�t�9��D���H�缬ʶ�?������f�$fG��;%�ߋ�s��AP�X�>m��7�O,@y�\f�LT�z1�~�J�R7쭹�Z��7�iO�:VL�q�=&�V�Z�ȩ�6�������\��Qi��4qD�(�i��]�5�TZ����&<*����p�(������i���o0�ϥy��L�kA\6�7>b�(	�sm7n�y�x-�k�dr9��eRo�y�\n1���e��^�{!�Z~b���`$�z�Q���=����!��	J�39�(<�̪���DA:�x�
�2�ˣ�뭟�&|=8X���&X�P[�̣�*Ab54��o�pF8�i&��ɐV�ۚ*-�U�:���,^r�\r��B	[�n���"�X�o��2��IEK�A��<S~���8�LQ��F/s.�ϐmFmyeV
o�Mq�.-MT����h�po=�������4��4�WI���$y���#��e���uw�ϊ�W�e�Wɳ�gڙo�%�39�~ߕ�u��yi���tߛ���㑠)����� F�슡�H=o�5F<���2mZ��Ws�t�N E������ �E{����h(̔g�6�}����G�f�J�m;*�����!��ұ�ee��u	�%�VU4̤y�2&ᮏ6]�ʫ��տ���|(���+�x�m�zM��U"�*��,����D��TM��U����Ri���t�^��!¼Ψ6r��tؑ�o��nA
;�'�yv�����@@��Z�'"#�%j�z����S�I m`U�W�qo�=�Ci�i��g�@��I@L�kF�w��v��D�8�$X�i
A�����Y:�{Bw�e�\�9Y��?�Z�@��HTL�7|�@���>�W��c-�����)W�p��s�;놟j��\)���ջe�Wg���S]���ܐ���|�Ն*��D�x��\m$^���e$g%��r'�J&S����}�G��-f�L�� �����5��S/�������[�|���H�=A 
�t%�9ңo�<�R-R��ڎjc��`d���P��¦����lr��i��$����q��85k?3�/aMO�'s�4���mWv����.M�6 ���~m����A�9��M��[{�=�&�s/F��~P���R��t^���p����|�e[e�~�HC�WSǐ�|U;;�~�����������x,����L���6�Al�Ji󒀯?����?uT<�ƃ488������УS��z����\�o�
%� �־F�����"D�d�k�ɝ��b��`m�H�0m(O�m��k,KC$4)O�`v]�a��r(q&UF�_��E=LH�`����в|����:���X� �|�tvp�IY��9���e�`�s���d���5c���=��>���Y�G�'���vѯE�2i��>u��6�[&���`�F�3�4��c���,�Jf,����m��kwu��nd�L@�/2�hm�wk�U���t���%����;�bm57h��S�LX��2M"�^���Zˇ+n4��d�
�~�_2��1=���Id¨$��V��s�(��0I�Vc����PG{��EQ��{d�E���ɵ�sd�8���7�?~,�
[�
��/|�J xϹ��}�Ȅ��0}� f�u�(^�v�d��#QW�K�$�F^�WI���Z���=��DGG�z6a],��*wTٸ+V:���ABf��T::4���f�|��c�!ZĹ�E��X�b�(�Վ���rf������y_)O|��_Bqr��;��d��b��dC�jMD=:{�a�|��q���.���)��4n��=��wSm�
F""7$`/
��.=G@��pR�e�QV���o�:D�q�/��Uh�ZQB����Y':/��OJ�៽r�<J���#y7�x���X3��Nÿ�!?�T`����@�iڵ��>xB���2�l;$_7��蘜�+Ú�����ˬ�͉�E���\0)6�³�ўD]��{����]�J˥Dn<$���W����)�Q��G н�1���Z�g@�k���q�Apr�`���\"�B=WUt� �ұ��\���
p�/	��-t=����00�aA�h��d�C�գWe�Pݕ�������5J������Dw�B��a�\2��Ot������f^  ������4�k=��,9o���a@�4s3RN�T��4R'X��3�>��Ǣ���aUY��<���F������+U��C�׿	6�8���m���.C���k$�b4YS���z�
���lDo���x�6Ҭb�	 L1�f����A�^4�
��T�ګmo	���|��=�⩗5�曱^Ӌ�k�����i�`���kn��>��Ik kͩJ/Ik&�;���xU���"��,�n�;PQ}ى8��
Q�)$��}"��	.�|��i�v*(A[Nĕy�U�	F��h�n~�n.s����S�g���X��rFƽ?��3�A�&���E�v,������%�'j�W@?q{v�+�9�:�����H��kL�ރ����6cu�#���뚦	�-����˧��)t�t.���*��)O��$gbB�Z��=Lc�P`�-�{Π�eK��Ɉ�q���y��
zt]M��%��0��4��v� E��� �['�?��O�%v�]<4V]F>�ί���Ao�֕F%ļ�2AߝkͰ�lvf�.OY�:�퐾$�/���|{v���|�>[�$MWߑ��Q^��8X�/R7oMza?\�0р`�qXl�@�r���)j~*ޫe5ls��c{&��6��`���Zn��mmv&X���7S"'O��G��--����Y'��feԶ�ҍ(.aG��+���5��r&�8\�B\|A]��p9�j�5z��9��P�m:��TG8Z�J:Գ�n��m���Lr%ٝ!*�F���$��`Jx�ʲ�|�U��Qؾ툔y�m����]Uz���|��P�'0F@�u�kA�������Z@�<��{|Q����uJnJ�y��	��� G�D1�9�O0H��)����wK�0B�8h���O+���4'jD�W\A�'�ms��zeC��+TjB�K�:Ҁ��VY2�!9(c���ɤ���e�������+��P2���A��u�� �.e�G��Nw�\�f��s���(#*_PF&Z��1l��=G_x����q�B�{���ǤW�H�k��bY���Err\6�N:YZ�E5�330>|o{��r�s�ʀ�zz�<�eD��L�K�^|R�����F�TT!Ev��`�n7���4�Iޚǩn����{ڰ�;7�,n%����4�v7d�*|]r����$�6��_��*L�}��.�q4����E�9~�^.�x`%hj�eAB�(��{;'ڵu��R��KFL���T��}�(�4���J�3/�7���Z���w�����o��-�=��@p��� R��hW�y4{S' ��T�D����1t���?q��T�eg�������X�8[���E�c�ʫ��J���Ȇ��p�0������ٟ��3�L����5�KC�s��oq�����U�x���ƾ�/"��-���P��bᝪ����b�zrF-@�����z;����cvAlH��J�>��T�nng\��o�`�?;�'Qwv���% sD��9��byҦzL�u'�L�Ũ:�4�=ڀA��7T)���r�e�W�$<�D[)϶��jð��xL�6���n�j8:wp���ϛ�'y��}�h��_����+\�}�B�ՊCBIߊ#f)���*WQ��	�Z���G�/���?�R� �h8Z��Cwj_0��Y�� e�l��M�R],WMvH@R;�j�g�6g�3U�V��2���	� �I+<�4����@�Be"[I�l�)@`���t��$��}�+��=���   �����Vwi�.�΍��P� @�qQ<�q�ϧ���L��Pg���G�,��Q}�?+sY?"�x�s|��O��l����ƭMj�_h�x����H8�#�}J�ez�0Iᇫ�cR�Z�8Bų�=_��w�cm�����=&�*���p0#�O��}���[C����Jʖ��bb6�b�D�xVM ɷ�&r_ֹ����(��a����([ֻ���83o;�
�Y�]a�F��_S�gW��]\S�=̍?���-M\�F��qs�e�M�����#�G�'���ɬ��{�Br��(L�m�n�|�|
�7n����x��p?&K����7��M����'+/��Vń(z�|�,�l���9!�r����@Gr���1r�;�,ݺ��{}(�Q�6l;�_�
�x�d�Y���m:X$4�\)��3�j��r���y���9f������������� ���(0�`�Տ4�f��1���l��U<��%�S!������.�^�+sU���%�&"�C�>�<:�Fs }J,�'R{�lT��Ah4�O��J�Z��W��Hx�O2�6��خ����KZcگ%��U]v��}���T��q�{���	p����"�9#���]0���4]�J� i�h.�����(a���f�.{:	��9P�L���s�6t��`55�I�O�C&�u�.�}B^N��xy~�J�t���(G��-���6���b1��YL�nV�%�a���t;&a�f㌥"�~N��%�2Lv+1�[PF�<�a�'��5���"f�w���k,�HI���tk7�{���&e�>���8�D�k��Th�]�p	�?��
%��<~cI������=	v��ai���v�0�/.<}w���9G
:�wF�Z���~�rt0_��ޢ�*�)�
�[w��2�F���ו���ve`����7�gy���ID��!��g�`���=o*'��?wr(5½��m�՜a�S���.�C�i�x�
g��,.f������SU�<��)k�,Br�%�N\�
F��FfB�F�h�T��~��g�;���E��gb�tuE�]LK�HfA˨*�b����I�5��/��ʼZ4�z^d�p~�MeS���L�cw��U��CՍ�E
�9u����r�%�n(�\�p.4{0�B��:��P<��1%�S���l��Oq#��J��L�ZB�L������t�ɹ�N���;3;|��IуU�}Qw���������߮�����u*C�7:N_�_`:��+����1a��[	�i�O����#Q��v�0/��Uۀ~�P�w:���$q�p��u�!'T�'�l�p �0-<�mO^��F#�1���Z�Q�e���'�Uc�϶�D���).4��yZ�X��l����*"��wJ!�=V�ŨؒQ �[�0Q�;CD&k�����ѩ;��r�'�c�o�x�n��){.�2M�RD�����v��
m���s�$~��J�6^z���-��������s��@٣�".�!ʕ �w��j$�۟���.\�?N������72Jh�.b���7��<!�]�|�I������@��E~iD�� =�\�㯟;6����o� sb"pUcG(�IİTG���V�<E�s���Y̳:���fu��2!�n���H솨Hv����ATP�������_�p�]���J';P!�l�}�E��z��1�'��IDb�>M��2�� �X]�o7�-�&Ra�W�9�]E��z��{�K�F�N�v��Å�(Dpz/��O~�K�))�{��8r��'��Pل��ؒxh�v ���n=F�>=֑�[��x���%���[ֈC�>��@��,�j<�u$�s*�O�+��1��$㤵2��<)�Y����� O�/�._mNU����1K�Y�2�U�<M����)�4�s�y�����:���4�RcN�NO�DGu�c�_�_؃�F��?U�l��?,\���1��bx��it�&�`>��2W��
��|?�`���%+#B!�R�(��_��yb�'�`t2^C`NGr����	��lM���z[M'��V�h��{�O� �M��ʫ�YV����]U�j�J;2�ղ�'��y�-Ų�uލ���sYE�<E%\t��WNeQwY߄��τ^{~2�Z"����u.�"(aB�ˀBOs[�����-OqNx]���<�wH/��B����o^�~A�s��Ԛ?�Y��G����E���S���C���]Zg��{��0����ؙ$����B7��#m�V�����@�8\���L��ۆY0%g7VT���;�$6�~҄��H����	�6�['oE�:6�<B�� h0�#;fo�o��>3
\.Xa�UM� ��@�JV�@���� ������+�o��{b�])ٙ�X��JUT)�Y U� �r%��̋�,U)�cei��m#��[�rer�6�!0��p|��l�D�]&=�{�8���RVє�C�����|����^CS�c�R3:��S�5�͇3OpT�o�(�� �:P[R��*J����8,�؋�e��+f���ORS�M�Z3���Љ��M6F_��� u��8��@RG�1�	X�"t]2=�#��q76�L��#��<�k))9a�'��*s����e��*����fO�6�|�0ۏV[���x����n�v.��F�jo�i�z���W�S=��~�P-:U��u_���Q���j�BFǹ�9�r������60�����tM���,���8iϦH��"�$+�H�rw����8���@�����RM���/6;լWFM)ؿk����ΰT�>�u1�^fU���y��m�b���i%����D�rY}��ul�6���~�@�Ň(nVn����s�xKi�]�Y��%��w�Tw����/���\3������V>隵X���
u�.j
���R���v~9VF��XΗ3� ��{�854���Mm��_1w°+����j��"2����d*�ð���D7	�70x�e/�O�%���.��N���pQCb�������ۭ�3w��T,�s�C�sC�����d�������KmD;�8�5�o<�}��:h�W)�<x?��{�5I���^G���e�����͡a�j3�8 +��K��V4��i�!�2I{�R� ��/9[�%O/�ʧ�{j�_zkJo$��s�l%�;ʾ�S��J��� GR���8���c�H�r�=i
Kt|ƿ�-{�3v���I}ƍ�0��r�O���G��tG���]�7��p�UH�̞/�߂�1Aq�a�Z@���V4��O	�/%�@ [��~[�������3����m���G�SW��0U�g� ���[����L�3��3,��x�z
з�\�xܢV1ާ6ɳJ���`�Ÿ(�e]e���\ZY�������M�+iU{F%�~~P�R�^��ɿA��zPR�������V�0b��c�6|��Bq]o��G*�� ʝc�}�qG%l��9Z�����b��2=�]|_t��}3�Aݬ�sU�(����j��h������t�5rȯa Px�z"E�6` ����'x���Dd�+"�Q��*y	]T��Ϝ�ێiO�Q�Y���0�R�.��,���>��|�~ڐ�Ra70��D�2���f�����������!�aO��W��F�d_�h�j��LLCl�V��c��c6Ԥ��h��,7�>�
�#�/�����e���c��n&B���\�א��� �+ϙ ��ǝ���1#+�N�X�8�R!�՗����[�`d�"���%ȴ�%%�+����5�>'=ƀ),+e�ǻ������e�	� �j�ḿ��c�@����	f|g�H�@�;����y��^�/	�p��
�Dz�5 �9��d��2Om Xm5���,��<��J�"^�L<j�j�o��@�kt*9��k��K����N�s:|���Nت�g+���}����H�U*ޭb�����u�f���5F���F�[��y�-=�����/����ڏ������v��W��
���d���.W学r��h���
�~���-�(�E|;������cPר�����!fl�ߕކ��e�'�9+ � uҝqQ�����Mgs��m��$����5`O���#���G��D�O����9�ꄚ�W'UK&��Յ����r?��[S�2[�%�A6����'*�|�fg��?v��?;�su�(��|o�ƪ�#����;H�,�j[!m�H֏��7C纅��e}����T�j�Dqhe(?��Dʮ����	p���x�r_�$���s��庇�J��"�!���+{Of��b��_�o�ѷt��M&�@b���hD�_��ӹ�~:��%V8��{eg�I�u�a�:-��[���\	.��]?������y N�9�\�Qg^ƑD��L��iD`�g�N�<��>aD�Ԩo�:m(�eCX����P$��2�OCK�L@߰��G��ڷx�Z��ۘ�d��,���:'J+vƖ��ǖ�C�K��	�="E��%L�˗�A���'u�c�,��=ǱBB��k�Э2��a-�hu$g��)|/놑�>$j�Q90��d6׎�Ȳ�SҴ	ܑn�5����q��L�P�Mr�=�90�}G��2�����9*$���^��)~�����	��m��}LS_[��:G���B5^��;	���6���Ҋr����2��m>�a��7�ږEK��3EuG�������{����%\-�Q��Ɨ"��L��n���+������.��`Q|>�Q�zm>���R
8N�vϦX��VN�[m9;�O�|���92���?4<�c����\��P�:-�i ��f������3\Q����@���т�7����W���mTZ|���X�`/6��dބ;�>�CD���
4�5�(Q���"d�>�f����� �p���[e&	�E��HrS@������3� ���Ĥu�@�j̕\iȸ�-�WZĳ�h&DC������&>����P�7�:r����̼�*b���iƭ�� �-���W��e�d�^W#����,3�g�����O:�4��Ѕf�"�@�J��'!ٻ7RSl���y����QY���I��d{]��螢�)��>xq�3I�z{(��>���O<�X&�mJ�Pԣ�;������W��cs� {.���/����c�3۬�����{a��v�2���s�H�%wz��������^�>�*�ѷ����W9P[V '�i1�b 0� �>l��2(E޸
o��U������������n��{Y$.�P���k�?3
C�$��T.>Ș�8O9��-�c@��#��p�ɩf[�p���Q?�'p+��F��hf�H.d�n�.}i��Z�O��|��@�X��� 3Z�ѧc^�n����\�L<Xy�x��槮5�,�4�oٰH�������Tw�s�����C|��út9�-�ű�p������ծv��X�%������"+�t���$J�rZ���%J��Yʋ��Y�77�ES�̬:�X�`zE��?�(_��&�?��5��#ࣖ42S����R ���n,1��M����<%��ԏ��W��85P�i�i���gk��rXx�C�H��D��NBİ��NnOP)-6��E.k���~�G���L}�'�o>��� ��&�.ꬆ��<��b�SЍ���	�[�����֌��mO�NS���)��J��움��)�q���$E�w.�߈n����&����$sTY�θ�� WL����Z���jf�]E�@,M�X�[�-�;]>�2 �3i�lAl�m���=.��\��sH�� ��?��U:,�h[J����Zrꀃ%���*t�:B��%�{���t��X ����y����s��Z1�:�Ӽ/�*3t�s-��	T�p����nL��<�6���_�o�`{k�zQ�|��V�n�@�T��P�=�[X<i�$����g* �ls)6��K��љ����ڀ�׽��D���u ��2���H�枕�!8!,	��ޱ�Ǟz_3`�5�[��.�R�8����K��3�#>
ܗ��3�rI'�%�+2������Dԡ�������+brZ�٫������i���aX���H�h6�{�ؔ=vىx�� ��FǕH�?V��{w\��]ť����{VN!c�Tmf�+]��&� �2��IG�d�9��+���/�*�`8��ˬ���ܮ�%w��� q��U��Q7�r~�X95.XuGH�8ۛ�{ίC���LSɯ~�M��(Fy���P���du��*MW��gox|FC1͉S9�DxbH�6����@D�=�o�`}p�eGaD�^z|D�c�qJ罋3�o�M��'�����EP�G������I�"��/L�H0�z��}Q諤"�I����������
1���!q�.2��M�-<ޛ��kW
��G��4(�(�
ڙ�J�?�7>v�r�Z�֙��sy�J���`��_���v������|G�mʳ�,󝊡�(S�$�ôI
3`6j��dm3^����ޮ�Ȏ:�^��Q��Y��Hѿ~cMX�N}C\āuM1��~�利	 �K>�@!��}{�>q�6:�~h^F*�������Oc������]
Ѽ|ަJav�U4���D��rtMS
���4K���3��b/�y�B����������)u��8Y�������f�-C����NS�7�����&�x�WD�@Y`�4�8;�H5^)3l�ō���q�@�Z,���Q���G4:^0��1"�^��6��a̋�,��R0 �b�b	� ��	ԙE� �R��m�j��d��<�z��jl�L_h`�&��ǁ�vUO���H&4QV�KV�I\���>��v��w���*1R��i��+7�� :g��R�[�̈����9M�6��DUXu�+��gKq��33§�°V	�����	۬߰���B���W�4�;!7�l�9^�Wߪ��Vz��"�j�F�I������\'(q.��|�|�]H�uw�!��� ��-g}�u���9?�y�hn���/P7������T� ��2�a���� �)�ȓB%ٍ�yi��pR�����*��'��֣��T���򳻌���w���!�����RS���Z�8N~�F��t��khm3kf�[�i96������1�<e�ca���6�-nbI)oqu�%%V=A��¶���&�S��"^) B�Τ�6yBN(�_#���4��M|�8?QNe��m�(�\�0�<�dE[ڬÂ+�C4��r�& `<�6���f   ��9ź}�vB��ѠF(����p9*f��"v��?rk��h�}��✢�\���$o8�O��Ӓ��4uO��z�h��Lװ�Bb����ͲP��
���
�,1t<Ym\_眶�c��e��;�v�b��`�s��~�+����j2F�h�a dqLIl�v�4����/�R�`T��JV�j̾��@��龳ީ�Qi�H��R�+yO�uje��;�� |e ��ˊo�&��&l^x�C����`j���j��������|j �-Y���.�sm��}T���D���i ��¶���B���]r��� �P�ښ7��g�:?�2�Ӟg�}�����Ҹ��z^��Jמ�?��7z�`:a����_M��e�I2�W-6ʯo@�)w�/V-��--#:�[��UP���")� ��%�V�e/�PN�FOg(L�>4�ud�C��b��E�$�q��=��S�ʰ�D�j�O�8�4�+^
PI��� �b�����)�I�p��Z"�l�-�.�}`�Y��/����kO�ڰ2�7R��ez�Y�֔p&��c݀���8Ō��.z� ���]�j��v�
��+�zIz#-vp�'�g�G=�����v&��#
ր-Ԑ�֨؂$�/�ٹ|��(v����\` �0ꗖa�c}�]"?.��Ghv��C]{&��%�u)�a�E����[�ZX���)Ps���Q7�!<T�a5K�]wg�j�l�t�=��Kr��ܫ)RX�ꏎ��`z���p
s��J=ی�+	��7����6���5��Ç�d\�� B���ˍY2�Ћ��F���i@t0}���no�R�ͫwO�������W�Qyn�V��U��d]F�����S�
%ж2��p���x��QsHˣf�UV���&�rJ��s�Ü�9X�r���|t�m�w�.�Ў�g�B�+5�H�׼\�A��_�X��^����䆆�H�2|�x�>n�?n�Y�G:�ݖG��YI�x`�~O����u09G��\��zJ`��j��fK�РY���I��7��r��A�1� �DV��A�e��2�