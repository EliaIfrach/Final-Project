��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S�OO�$����d}�嘩qw��J�����j9�ܔ޴k^v^�����I�K;���\|�_X�`Z�3;Z���TN���P��,� �A[�g���k�ȱ�C��2�������5[43.��Lw��)@Q���%��C�9/�ǁ��oj,�̊1哫쇏�K]r?�GKV�b��d��N4-MNy��g|qd�j:;B�'���'l�+�B�ĵH��]���aҧG�!����Ӑ�3
�9���O�DCTB�6�t�9Hpu�l����#��p�����D�\���8Z�p:��7Z3B�ȖICǅ�S�~������˺ʴͦ�O,������;[ڳ1�Ui�W4�$o�ꊪRĭ*m?�69ӳh�W�6�`[H��cn�ڸ�:Y�+���fT��֕Tb'����z���㨂%EC��VM�kK(Q�cϴ��	����n:�\vvnS�&�-b�YTڝ�&���C�p5>HH����e���b���d��JoZK_��"ox9j���n1|$�b|��)b����D;0�!�%� 0��=���F�=��@IR��Q2�^�i���1X�NK7��t<t�8g���]��HŜ�2.w��6(.�� 6��K�i�y�_���2T���43�f w��
��B:�qjG�y�V�o��AvQ�3���,Z�t�j]m	a���9[�9���ol��`q� L�t�q�j�Y����a���^t������g
�`���em�QQ�?*�;��_�~��7� ��m�­��;C�c�+��N�����	��z�oS#��76�:}r�e���t���V���n�eMQk�Ȍ�59E�������Wg�V�&R��	є�Z!p�B�kA �tttN  ?~8�1�����K��ӹ�ܫ\���l�����G���׿�OBóM�(0�kJe������A�{��&�~��Qუ_����f>�%}o��~�w���}&c��^���fP��,fA�!�x������������C���W�����[� �^]~q�
b'4A��Lg���	�8k��L�T���l�i�˸+���ud�׹Y�G�L�/B��>����C�$8+�p�3n>Ih��v�̽��c>���1����J��������EC2tK�����&
a�y>y�k3�pg9�$#�m���?d�)7�1��2�1C�h52���Msi�zB�!z}�/��s1�W���êd�)�K��D*�e�eZ���TY�T�Z�-�1�p|�I�?�n�����a��]N��ݤ�A�j�,}c�����C�!z�3w��`��� v$Mct�µ<�d�D����!%-1IEZ��_�K(��@_���1j)�[��ͽ,J�컱n���M�^��q�51��Q@Н1�^Qӿ��`���N��%*W�k��a���.V8`�ˋ4c&<�!{,YNKO���:84����n@~ks&�&��-]�>���V���S��I�䜀�5+.u��|��"��]�"���u��a���h9L���G+_l��Z	IwT�*�ݽ��.\��!�JA̺�o|Y��̄<�0ը
�W@G��i�i��HP�؛G;����K�S��f�F�I�J��(k��k-��K&��P�г?��������`�)�5��#v����#wЅ��\�̨ߜ)n�^F�Ư�ga��Ū���(� v���!���{� C����Me,.^p*W�O�aL��x���$��R+1��� �t�x���6g�Z��O��|����L ֕[YI����7,w���1Eq�)�8J�p���h{'��u�Je����fY�­�V��d�	D��RC��`��l����cM�}�i��Y޿�)�X�	K����u���\AA ߸�7<g6;Uؽ�l=��>2��;䃬�n��5��V'%S ��\�}�_���Yʃ|N���h-g�
kT��c�>֡�H�B�.�+��<o��k5���.6q�à8�3��@m�?Q�<;�Ӥ�E�;�}i�i��{O� �6���'W��Z��͝�����zg��(@3o/Q��Ny�J2\�51w]a�z,�Z_�cw�^r�n�W>��5qw(�����f�i��d�����M�	{� �Y��jrtq�Y��n�k��)��]�9[�~�Z~����$��O�)�r�@���!~Y�%�|��Bx}X'�!��s>�*{�Q\耴�w�W*���0o�_C��[=��CS�Y�(�Te��k�2�~{t}�E���N7�'c-�7Ӽ~��H5����S��l|/��Ӥ��rM�����cwRJ���%ɱ�Ğd9��Z�7�ڰ��,	����8�I�	*1���(x�0��M�9^s��؊@&$��[��Rp�0���9m��/ȁ)(��?�aHJ�7	�Fb�8�;x�J�������s��OC�����ixCD�2�9��_�S�~t�r��֕"{�^��>/�l�6��6������{3|�����p�?P�
��:���<ba�o�7Q�?mG� ��?��<�he '��Z�/��d%���6�L�Tx)�̱;����I�u�]c|���">�w��}E�9J+$Z+ ���F��n��3	���i���u�6��Ƚ/>��K[�6��7�
V {kW�&x7�������[�^���(����/U�bfE$���ԧ0��\9��@S
��	�
�!Mg�����	D��Ӗ.*P[,�V�˄9��̔�M.
>�^>8�����4䆛T'�	1�W���՝|0XM����[0��4|�f�.��4V�������;����Ɔ?��]�J��|�Ǐ��¤�J͠O�EZVZ͠b�<�NE�YB� �/���:2T�����&J��RܶS�߱�Br0y���R���GV��FG�����2�8_�Q�yM,��E���ށ�4;]@� Y�� ()a�:�2E��̓� մ��z�m�̫�lk�V���'I��i��!B�C�s8�s2�_00�vyV��$8WB�uɁ��RuΪ������R��X0��S�G_�.�hH;��&���{�H1��wFL#�4�K��Zp<y���O��N���o��l*(���dZ����iB�}�U?�_N@^�6���{���R�Qی(o�C"�*g�g6;��y���.�����;�W��.D۟X�M}�ڨ�F�	 )2�W~���)�β�檔l�YU��$;�Aaj$�|,�U Mg#p}����K�Q:ހ��Ҕ�I�9<z�{�
��K�҄�WD����	F"�<(U	�-´�S��t��)�?�AT4�,Tl��䭥#���4d�>� �X�������y�ʺ��a��Ȫ����Wc��<zմ!���'+�(N�������*�������W�7�n�oWͮ�h���$���b���v��Z]�u�~ݶ�*$�W�m5�&�G��K�uc!З�����2��y_8�ZXe��㳴X�?F=IQ\�wP&��S�<��7��[ZU�"���n�	���&d��IS�h���cBAKgr�a��n�vL�������:^�R�Kut0�W/,j���7^�H����}�,G���:X�x�o�²�ul̱��#��r�d�{Y���ᄽ��,�c�҆�ٰ3"�Ҽ�
 af�n(��Ȯ2iS	���o�T�)`p�Ri�@"���Ō�������?�'��t6'�XKf��:�1�a΃ow���Oy����]��Z|h%�V$B�T�]6��e֒�[�¦���?��D��ܜ|�R�<E"�Q��:����\�!J;`�B|Z�MA��<,��z�q�9�R��6��;�^ҵ�n�,�໣k�  ����b�M#����_�$�����ʞ@hX�{��v�M�^�-�bo�`���Ǻu�����Am+���,^7ʛ)�,{�;Ӆc���{�����w����p�K���/S�9�7��=��5>jNN���a����k02kGL���ۊC�3���Ƶ�<�m.�iA�F
Z&��@�˷,�.j����v�?��V�����X��5 t!������KՄ�����ܟG���o�&;��ʽ7zJ��x�J�F)�k��6����G�OΪ	eF���l3�-k>���IR���"�=�NC
`:g���<�['��U2AX.��>H�U'��m<�����|��R�����4��4iq�\+.AK�d�(u��,���b�	̈e�ɔ�3x�ũj�.H�$�$�r��"���)K2�X����i��e�H�4Jw$��'�h/+��!;@)�9*U��j"܃�X�wK�\� 	��M��M���E��koZY��6=����<�����T�])��z���c��V�n���y����OQخ\^>/.yN��y3jWd6gU�}�W:�2ҵ
��[�j`�ǂ���?ܧe�	��K������W��[�1J6��_����)��<�,D!��+�瑥6 �[�?�l�u�S�#jz�a�͸��r�gԾ�� �q�*��!���Y8+��$��fEEt�]�MΧw���6A&N�����?��v◔eC��'�]0B� 낊i����jDI_��S�����5�ϻ^᫴�t�?��n���?���[Ch/f���dwF3o�E�!�z�=�xd�x���J@<�C��Ӥ�A�[
��q� ��x�ĩ��ʧtÕ�A����ʧ֜��sh��5�c����5���:eљ㼟	�!���J���fpg�]�� I���,��ネ>6g�E���ӌ&[:U���a�te������$�'�V�����~Η�Բ�#�]���7���<��1�� �>��oɞ�XM���;�?%O���_(�'�����-{��U�'��iT�u���|rD�P!��C�U�K�y�����A���ڻ̌i!�/*��7?	��&>�Ӡ �#+������bǌ"�����i�VN䱝���ш���d�8q|��)���R�Fq<�k{p����B�������҃&���V�2����;صR��^p�ʶ.��u�ZQ�[#ٴ��E�����xŅl�9�N^8��ґS�(Nz��k7�� �d�f�h:��y._C�73��k�h��3$3�}(i3�����س4%c�p���][�����R�.��R,>X_���Pz�;g��5��ښ�FɖhAQ��:o����Z�7�u����D��nCw��<��?dD�k*6�hF��C7UT��/���>^�B��Y{Ju26�U����h���i��v�B�ݧ�v��% ��6m��?4ih�a�� r���B��ʜ�GK�m2+��"���4ؾ��[�� Jb��_gT�e�>�a��Q3p�v-�-I��x�m�w9��]S�JU ����₞�F��3|�����|��ڮ�`K�j�0���䐩�!X	$C��ܹT�V�X���3���z��@��F���t�o��ސj�>�����B��]���D*a�X~d��� �"�|n��(�8 B\���ߍ�$����<ٽ
JB�%��>R.��5F�e�c���O��r�!@h{�ݨ_V�V��^|@�ʤ�/�~/�&��ߟIR2x�pw�~ �,�QA`�E��-�^d�|�8*�U���+G���Kf��B�������q�-'���7���J
��a}��!��k-=�a�ֽ�}U�o�ˎ��7@��&1D���(����2L���]�Z��c���[P��p�*2x��kr��2Ϧ�<�a��� !6r#zl:�/�b��7���w�l��+�EC0|ּڪ<�A�`�\^24����"��b�b�{|���l�L��G���T�? W/N�߼�%��~+!�?�� by��e$pkt1s�>�&d�Ʉ�+�S�)����:l,^�#�rT�7Q���-�v��V��9-
>y���6�:�}�Zs���O�jh �|O�����擧��=?o���jB��bv� 4�|���
�-v��"��K�41�2��Z��C�\�7�;�/^Ko7ڳ���$�T�"C��\�E�!�؎���*B��".�L�� ���u6l<T8�`���n�x��v�N��@$�N��Z�&+�()�;��pu,��
 ^�L��#�Z����ӵً4���^!)�m��U<�)�W����b_2L�B$����@��Q��.
�Ae�x�'�h����Y4S~��I�G�.9H��G��J;�A�C�И�BW�f��\hsqJXk�<$MCIL�JOH��T nkG��|�����x�+~3����(ځ���r�#���_�p�q���@ӶPf��_8�����(�#��b	7����:.�L�#R�s���ƌ����S�t֦���^�
]T��:ES�c�ڇA�/̲�^_ِ~�ݲ�T|.�hح5kO	ԘϏ�.@eV|zO��gO��=�U�i0��K���&Tg�Z�|e��֬�~dy1HOe3��OUf��o{�wQ:��y(k�̺2��U�B�������$fˎ'd���/@$�9�fh20�~���!~>�0$\G��4Bv.�vj�fev�
��C�f�w��Iq�::����I`�P��N�^�j�m�[B�Ooߍ4o����;��M|��WO�"��JY?j4�&6�������iڀ�i˖����[����㹦�Z��iT�
v�T}�A�%������zG'��
n��p�
Z]P[yEW�G
���*P%1�fg��j_TƋ��3���W@"�-v�i'tK]g�Z7��\S� ���{�c6s�z����1D���Z@�ڛ\�3N|�)t&HY���t�A��g�h6��`���<m����#l�7�y���~1 t�]����b8_.g2Q��i�2@�M	�k���P��A@7�bu��n�.�k�sv��;�-3"qA(�H >����";u��C�g��52�%�jA}@�zu��ɤ:�����}��=�l��Jg �ҧ&�h�;~l��l�D��vW���(z>|g�p�i�TVȗ��Y[Xa���( �
�&�'���c?�t�����mL�no_����Х��S�e�S�� �)?�S/��CHC�����H�ˊ��q�lhC��v�`;������y-�¹RĊ�g��J%B1�Yՠ�o#kyL���R[}���e{���w�rL�[��-G�b&��w+S�6�� ���	�+��
�Ig�N��[=ۤ���i=P��M���y4���\p4�|56�6�SJ�ƫ?W�bF��:c�n~���pN���K�#�;�j͒Rw3pO,n�}Xʏ��w�xi�Xs�;�V����͡�~�~�������L�gH�qL��	�t 6���f�]2vIx2)B��j����G����`��'��Z�ko˸^���o�j��Y���'c|t��5~k)���mT
���u��1kIJa
�`��!T�3�}G�~�Y��,b�y���#��R�~����,3���~~h>|�;=�$f\:P���l˕a��k��Q8''�R$�t��ܧ����u
�0Zn���.Kd"Kc�Us��o�'\I���[�J�i1:B��i�C��|��l,�s�[}TC�ͽ��l_S�AX:2p��,T�"����Rviͽ�9wX2A���>�y����D��	�U��tr뼶 �e�Y��r��4QEq����ѥ)�0�8/������&��V,�n�h�[��m���na��z�v�d4:�2~�_�y�
�HGG���k}�Z@��I>!{Ęz4�y�.y�>��+l�O_Ks�m��28��_���;�A�`]�|hJ#��i�V����Ph�þ����K���:Bx�.�]KX��6����F?��	�8�;9)����!�k���>�tS+�Ϊ��������	��8�e� �K��O�CPny�LxS�"�{�i����(�D�><T�û&c0�C�V����	|����nB,_�@*��;���gU��(�׆&��-������T�Fb
T.Ԇu��C�;��ʝS �_�@E�9���NA�rٝ)��؄�It#�f�,���>S��/�ڏ�D��س	�!�C��k1��^'�x+��;b��~�W��ݓ�Oj����UB9���xp�DM�����WX�b�Vf�Z~B/:���Q�k/�2{����셍� fCn��x��Ab�\Q��{/�Km�!��K Δ@��k�w���H'�5�`�K9� *�%�>��֯��]���נL~ԅ�#*�^���Y�c�Թ�4��D�
:���O
����PĊ�椘a��Y��ɠ���
�r�j
�T�E� ���0G���Na(l�=�25�����G�%��3@p�q_�=�����fc�?n��3�a�d�.-n�?�
C�Dì.�y9��%��Hu?��,$�p��C��=C�M�p�lj��-�+L�mn��j��E'D&?\�TG����=}�h�<ZP�Q���d���e�`����DҬ��D�R��z+1yq��Ũׁ7���`S�4c ����ط��	�����wĄ@!M:sY/�/��sQ�s�ǂ�����*�Ū��\lNz O���X�&�}��Y����T�3�w�WG�F�F�B��婃�­D<���I,�;\�j7�8D~`Z����w�H�t�e��~�E���o�L����b$؊q���b"�t+��;�>]�����{}���l`X���^�s�����D��X���w���f7��-Eїέ���6f�G2"nr_2 �S�$q!t-�ip�?j�d�FW��*(ь��8q"�y>B��̝ueĆgo��8f���E����5�����d���0Dc�b!�#$��y�>6��C!���7�>�ǿ���]Pb��9�|i�`�z4� �A��a��Iv�Q�q�4��uP�{+(����CM�79���le�~��tM����V�Qَ�D>r���*a�g�n�Ӑ�<O��I�M�Ohsԙ�kW�+�6�0�����O	��T-A�Sloʼ���S��}�i�s$5�&��)k�1�hkd�H�CY0�{���3gL��OCvjJ!�OE�H����:�d��k4��h1L�}�]��A�U�=:�?�z2#f���˕F;��@)�t-��)�T�Ε04wZ/�*��\[�#),��w�f��q'"n%��B�K-;��9G6|9�:P�� �1�����3��[[ac�{҉�9����|������K�dD�1������C��������dL 9�Xl�nׂq�K��E��g��g�*�+%�d[�$�\_��=4����.8f��k~V�ʘ�-鶕�%�Uӡ���4�a����)�z�[������$J)拝�h�9�̧LR��<J�,>g�}{5���v˧�x���$�6R����k?��v�G��z��]i)Bݩ�=����%9,~�����^�5.���&/w�j�T�D��rM�}�"��fS�������?�$����P��L|�_Ƹ�����ex�����Hn���˝b^pK�!�{�̲ɥ����,�Q4 Ai��7�x� V�����2�2�/U�m�����׏��K�d�k=,�����BA��j3Zo?U���F�)ț J8�c�{�^y?��Z����g���u�	at�V)��F�J���)��.�"-/b����*�i�/��P�� ��CY��I�ߣ;3�w6�t�O;�ʇ'��FDo}��ǶxЅx�FBKx��&FT���ɶY���H�p�W��r8!���n!5X;V@]#hL8�uR���a?5e�����Y�~Z�g�VW������%�q����gb��Ƨ?/����q����r���~��ϲ�D!�/q���B-E���}��Qôwpk^� ��Toe���\Ksuv�n�Tz�LM�H��>Iq���ş�KU0��@|U�v��`8 ����$�YL]�tĶ#R��"����:M�7)jTd;�9�U[�t˩��L]��r�Z�鏓9o?`�k\����Ҽ��w����҉��ʇw�������g�C*j�Q��x/泐²����_rL���T+B�ꭃ5�a�ft�p��(�'�9L��?�k���7��O�͞>�;ӹ��x[�%�u(��w��ȶ�*��/��}�ʋ+��k��C�����4�EG8/8�B#hX�kiCZ���ʯ�of�`���%�X}d@�^�?���e�V��]K�-Ϩ'����v�<�Y�읭���9���E��%�ি��A6���}���֮�t�T���P�����y旉S���{�5#g4���V��,Ꜿ�p�`	�I�S͋�QJ�+���e���{ԃ31�G�TG�����M:���9�=6��zJT���vR�|��� U��J������ vN�^���·}����!���B"�咵�i�a����$"��x������d��?��$	��Q���3�b�f�I���1��u��?�^gL�����b�h%���_u��CX\,�&	�(@{�!|Q5z�Ε]����6%\��@=;�I!c�����Z�4SGL�5����Jڦ2_���^�ܺ����{��U��t����Z-d�ޔ���4DG(��x����Z$�ZZCǖU��*@]�G�E�P�&��di�Y�B�fIvzȊ��f�f��R\�n�#ʪ��j���Gi����
��6�<"�de��C_��_
c,�a���1s%C��ec����h��S��n���M�C�5�����l�whMB;���O�²Lh+��U�Sb��"�b �*�jV��l\�/�O:����N�"�NԺ�蟛L�f�0����6�wu�քG�]�/,Nݕ��~?��w��_�.+����b���[����Ȃ~뜖���y0�ԏ.2zĪx_����n$�>�O�$��#�̅x�UBg��Z_z�y�]�x~��q�����nY�S��_������w�y�<+R3�<U�1�����R�P�Yr(�#�;{�o��W��NJE�9�s�n���]��ܺT�i���/���h�{�Y����GM�inU�p��g?����-�d&t�~����j��7�nq���m�S��Q\�m���y����p6&}�S1F��Nփ��������E~��	�d:�&Pz8Of�OM{
(�~ٓMh��\�C����c�߅<�.{��-�8A�w��c$���� nA�O�γ^�{#p�*KAڃ$'���mG�u ;��;��{�ű
ƫ��˕���
G%���.��{yw���w��]1B�1����1/%C��v[v#qPP� $Ok���i���F�n��?����6�*2$KQ�eX����e�`d�j*�e���	qN�9�n1���?�
.��#�j���B�[\���p�0�¶ԫԢݼO��1(|�Eat\s�~Ab'tK�٩��,I�P2��f;g�@��Y��Ĵ�٧��5W��
Q\3!��H�i���,�9�^4�3�9��p��=_���e�T���k�tЈ,��PR��dٕ�FyF5�rB�y�fnf}��l(�{y�S
u��Ú�LE���G�F��,>d��F*�#u
u�V��o3���L��a�4�Ak��M�O݁�c�O���\ٛ�73�X^o�v+�%ACqV�A��ڤ�c־|O}�0Wk�hÔ��',6냮I�>���5{��C�0yH�B���>�a,��X@ǎÜ�����->�u�����ʖ(#�����å�x���^��_��ֿ�v�� e�UT��~��D�ݮ���>�[�p�j.r��m��c �JN<|f<Q
1���j �D�g��R]��Z˴��0d���h���W�tq֗1��f*�+MM����~IG�0c^5��9"����G� ~2�d1	��*)5��21�t���T^c�i\����MK���L�0�{�am-�Q�\k�_ �0�5���<���N���W-]����\�ЧH&�)�
k<�䋃'�� G0N,B,9�@�E8
	x�\��C���Ӛ����R�T5�J����W���a�� ~��K����JƁ�7�g�~�SW%�>n�ڊ�;�ch,x�8�ޒ�,���.�Δ�eW��ӫA��C�q�=�6�/���<9E_��V#�H	}Et��\f�1x�<LK�6��A�^���m�C�l<�cK��d�yBз�Vt6���|a���;��n4�!������N~��י����e���G�)�)ۦ�F��Q]� ���6���Kn� �p!��3��Yi������`��� 4Op;�^h��ӽM�A���|��x
��ȃ�b�C��UVg0{~�D�����֢�H?��W���NY�gS��S��1����N�`h�*r�<�XL7Fۃ�l�5[�ܳ���|��i����A����j�՟���Po�(�,P�~&�5�u� ���u�F��,�7Tle�A`��
.��N���U��^oĠq�#�����"��<��e�i���V��f���:ߏ�Bfoql�E�3φ�Q}v\F%��K�np� �jSG��1BCyp�؛>���A�M�Jǣ����s������.7K��Ju�YyC���X��<.�7�o_���&��(�@�ד��¯L+�N���G^������V�<��P��e	�������Ļ��+���d��I�F�����[�E��nQ� OG
�}w4A7�J>z��w&��o�|un��]�C�I�$/�tV76���[b+��6u��@G0���������«
V���[�(&����O�Z��S��*^�u��B�J�-�49���O`i-~.���8p�2�;ڱ�D�L�G	�̸�����d"D1�~�k=X~�_�u
���z���N��@�s�����7���Q|���.^��8�Yړ�XYj����u��SU���qz��j��˫�*���2��N���a�����r�YxZ��^Ѥ�g�+���&h_܌�q���Ce�j-��4�@��Z������,-c�8o�VE��a�=�i�ա_�jr�4�"�Z�bdqK<�Ka�p}Nk]��&�aI����$��|j���Mx1iX��/����k�(���*�[��f
�`PG����ߟI�ݎ�����[M���xf�	�>��˺te=�!�r�	H��8&{IS�"����kdZۢ��-�dʕ������6T��嶬��X�\G����9�^�6ӫV�W&�̓�~�ܼQyFNV����Y;��Xe��O�)��6�l��r��0��mT�M�ϸ�7�f�Gi]A6Z��?���F��C�֗��ha/L�\�o��n�������mx�͢��W���{��ǖ@~4�����[A�D~*�,X�h*��iL7�Db��KG��`F�;��8�%#r�͡C��2HH �Y�{��-�L�@[ig V��q�Ge�,�-G�Dx�$���$�
vZ���O<��*��vK]M�l	Z�y���� ;�WC�ܪ��'4���y4h�榤�����^!.M�E���L�Ǯ^]c �?w�mD8�7�[�M��{��L��( eWmM3{�^��k��C�D������ ;�|�2�i戏Ĭ���
ż\�{sZ�j/�K�`ng���CTq�I}�1�����=�P]y���K�
���r�Q�!�U�tRyI�ps�B���M7>�HL;��<�ݷEd�*-�%��=ay���pw]��up^2�`4@Dju�"(iݻvsrc��5e�*�����O�u���+]��u�"^4��a�r`ҳu�#!���%�#�IK��'�L9s)��r^ �����ߩO�r4���O,5�W2j0���@����[��>M�'�<�!݂�;u��V_k?��y��w���F�qߏ�*&+pC��Vj�d;����Z�dS���]��O�l�+��F͞x@1��|?�(�3�Қ0bg�� }xD�,˸w�����(ϓ�ƅ��v�<��W�t���PƼ��PGP�՞ߛ�*��H��S��
�+C∩�/�V�`�y�q��j��b�Cc��0�*��ghr6��e��P�"V�����G+��*_���P��$_Ef~w�?/��@��f~��{"�5c� �������{xE�$\x�d�\��f~E �vc)GWg�P.Y�]i{��}���@��ߧ��z���p�r���ݷ~��p�J�I�1��+Lzј��lH�|~��\Լ��H����0��� �	RP!^vk�iA����svVR�Fo��[���|��Y���b�(�E�J�rJۚ�O�E��0LKY'U(��̎�*f��=��!�Tc*!�3�f��m�m��"ٱ�$�~�H�f�S�}�J0�%���O�@:�Mj������&��� ��>䮚K�3���#�gA
�"Tn�����?�MW�5�b�P���Fau7��
g� ��D�~�AZ~h>���fꯌ"=^��@��e?���=�p��dy�QRSc�c�\�%c�Z:�pFF�xz��]�gZ�P�m�<6zR��_���Z�F��˖�y��tq�,V�e
΃fܠt��p��lP޳��2��Wm1k荚�y~�(MP>�/9��b��f����{��D^�z~��ԕ���~�eEy��t��Ze�N���'K7�٬O;��B���n�����>,y�`nLvFϽ^9�&ɔG�b�끥��6�Y�A�3�������e,h��#̝�*⦬T;�OP�lu���zHI01��B\G0羄;9��s��A���Ԅ�Lc���?�V���\¡�Q"����l=�<��t�ރz�A6��8��h�̏]ȗ�ź�ƪ0Дs&QM+9��x�靚��kui�GQ����vG�6��l�Y��lX|�F���h��+�P,�z^%�{~_7R�z��3F�ױ::��G�2����	O��Aq�+h��.���^�``�ao��3}��^����:��{.�i[�z�����1��x�w���A8��ncBʫ��
Rǣ�6A�a׏�aT>恷�R���Ti�ǧ�)���w���r��tlX��d9(��4t_&��a�,�+�[Zɯ�J"�� �9�~�LI��f�	h>M|3e�y�ez��������wL�1`�u�[�8���6�D�Ť����r���:e4YĨ�)�I�}���R��~ݰ��C�4=t�p��Ѣ���T�}����lmZ,/�#!��;2NC���7r���c���{�|�aJ(����8-�DC}��r����e��<�t�`�����ţ��Ÿ؉��^�	r� ыL�]��>�n��q?��0I�-���}�ر��ؖG�T
.��{��%�܈�J3�43V�����*EE�JZ�@�JI���0��6?�ׄ����w5�<��$�Pj���U!����]],��Q��Qb����n���Zޜ=�4�00¹I_�A����l�<F��n��c?��,x�Y)��a:�Eo��