��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S�OO�$����d}�嘩q7� <���L���������w�Q��|�7*)⠠���Hf�(�Vӗ�����؏���M�(˔�Ywm���"jN^r�Wf�k���H+��M������}��GηF���L®������D�V�qd�kEMHA��
��[�H���+dKWJא������E��Q�]�B��_�WtLkg��MT�xrxC�������e��.��E�S[�!/�1���^A�,��Fu��8��E��N�s�|9�i [Ӿ�z0[���!������S�����O伖AGO�vJ�6�/��K��N�f��sr�:�W&ю���� ?3@�ۘ��c�*��}^}$� ڛ����c8�R�/��k)\�wӍ#X{��-H��QN¢#~ߦ�{�b��ۀwƆTZ�6Mj\U���b�,���|Y�O��}T����ru��Z1�w��E�{�����Niź��I��<��KӶ�M�8=���@B+��˗���w���-�V0��|����m:(2p����R�+�+�,XCRi�i�Y\���=ǞOp�V��%�qGO�/�Y,]�;�>�4�_�p�&�A�������=��m֗����Mu.�6�~>��W�	�TϷ�b{��-�=(�6�ud={f�T����0��� ��y>'�L�[�ɯѳ�oU��_-����6�!��&t}��Cr�,�e�_Hw�ܶp��`6�1�aLـ�����%dC}Y{yM�1&y���X����U:�ܲ�b�� �m%�S�gw���0�-�>��:tM\5�w�@׏I��CO�sW#��酅�u�G|�r�x�����a��,���ӧV!YɃ �*���-Q��BMaK�0N���P��ߣ+��B�ySGAѰ�9�$��F밚W��Sm��0'ӕG�C���bq'����@�	��GH�j ��(��]��e6&k��<(�nX�洛�R�:���{�ȍ�OK��)�➙/#��;)%~�"���/B��˖�W���3�7��5ϖ,�cm�6�O+�}�.��.��땰2I]9=�Qf�]�kǳ���#VD��8R�wQYA����'��RqR{�	
�@��PAXTE,�n١0�����|L���]���e���z7���밧n&���^6�qDÈ��p1f�m
�a��f)+8eܝ�b���ػ/$�7i� �ZIa����"�J���iy���w�&>��c�++ D�X�s2�'�(R�I�֠2浂�k2���Hw��\3����(\�Q���w�H�:��l�HG��,�b��*-�j���L�hx�=�/�Զm�Ni�|Oמ;��:)"C�g�(i�$����Q=*�!�R�Pua��y/���ri�E��Z{��Y��2��d��2�T�|��	�V�&C"�
���U˂�� lF?�Tj�X���!�Z�|�##w:��vƬ��b��������$e���~��vx9���|�]ꪭ\�����&/R�^qҦ)��/�h�F�!��	N�ؔdp#E�8
�ϟjT���=��m�[��$��Ry{ Kˀ�QQ��/Ώd"@ޅf��Fh�N�Z ����!n��$QB�J�]�'�>²�)��W�B���>�����R �N�
��GŻeֺq�(ff���<������� �T+�y�U2�OVG<��9�`J�Q���#Ϡ�����w��]���M�y��J:]lH�"�Pz�QTB����"i��y���[Ԡ34�ga�T�^3@����T�����/.�&8��{��2��QP/���1}�Ē�7�*A�w�()J:�g}
 ��˖%�}/�4 �?��I؀k*ާ��xcWm��l[k�{�mb�>B��/˘ <8(�U_�OfI_�ʇa����e�Ɖ��L��!�|�R��|sWA"��������H�z+��`�ŶH�PC���d9!o���������׉�;t?��+}���h����'b����hZ�6S�Q�/Q�i�,�\��S�r�_\U�A�s��q��zq���wG�;xY�I��/�5N6+��*�#�.�A�ֳ*SI/�Y�~��V�Lb�I�$����QDzU���hT�o�\�4Xx��/�
&��Ȗbo3<�L��I���-oe�B6�#���!�=М�D��`!J��S�n�B�4ߡUӸ�4�[q;f:M�`q���\a)���^�`�y��	 ��_LT�܉���o#�n�.[������x��</�T7"/��wSd .� Ӌ�)��wC,%mN��F �T��������؈<YVf|Ӭ}c�cJ]�8�`��3)/6��6���Q�W��ӭ���NԵ-��m>���p�)���m|vނJ��`t����mF��1/~;���'f����h&EhB�oZ���nܽ"��ٛ����#�?������R0z��{���SoZ����"*@� wM?���;�M�~�!Y`'UX1l/�4��&Z�����~+k���"j�ϦcF�+t��n����oe��f�G�� `a��p������=�[��9��t��K�j����R�;������$v�^3� m��E������O����m
�l���f]�H �}f�]	nF��lP�SSf��MH�Q�\���I�����}'�Ҕ}�5� 3�`��i�g�7H5��ԗ��6/�۝�z�T^�|��[2�[��'�oK"r'4�X�|��� �mM����da�� ���.��Z��L�)���;��{Lw�$%n���K�4�(9L~؇$b<��UZ??�p� y�{wG#����>d�W�;1��M��$�Y�N�����u"��6����4^[\�e/$`#�^�L�z~��٬��ުr?EUqex}	��Js>��A)�h�W�W�;Z&uQi ��o��8jnc&���/P�ѻ�u?�в���O�)**9��>�T�Kgl�@��W��ZXC/9�e~��/i��ZG�K��Q���%kE+��kع�5z��ϑi���M��&zn�?�u��fh�#H�, �u�@��h3����6N#F�K�v0��r�[�>XxU�?���=�ٻ�|��\#�*b4�a
D8,#��{��J%9��x���I�[$�ʬ���G��S^'H�E���čz#��s�H�,���4԰��	���&��OS~�9�a��嶷��� �}d�k���fW㥆��dZ����I/�M�p �����;��4~5�bn�;�;���a�@j�>�d��Z�dp%\5�������v�f�t�)$���lU���@(��P@�(�8"��%@to�Ka]`���B��n��f�o��%���D� ��Ցxlg��\� �B���]p5��h�Л<�$҇\��Y����%�������*K�3j�ٱ�7�?�m@ܙ�O��u���˴DR���8�]�{�a��Ks� ��X��4��^Uޓh��i9{i���P���5��i4�	�u��ԣ�I����O�G�6�)��<0���Y�C8#sI���o�rY`)̌��{:�$�r�W�cz�MZ&)���^����ލ����s;3,���a�����'�w�(��Y�oP�'RD��� �׵����K�
�)�?������Yci�z�lv��_�<��2���y��
=W��ݕ��x©r��'����=�c=$)9�@M����Wچb}8:M:�]�h˭}?��@.�'�(|�]��O����/�����k�GI��fbx������� z�
�C?}1<\�k6�.g��Y���=�C�|_]�\3����ɪ[�_uլΈ
/}@~�1��{���@�p(�SJ��~b���ppp7 |��q����(��X����Rf��B��[:��c]->tyw��._�Ü��:���k�s��zu����#���`��祄�~s,Z�H�w�'j����^y"�TWF�Xσ:���vv�k�K
i�ʣ���jߨ����a��@�tGvxr�??�,��a�*�ڊ��,3���Xa���A��q�X=&����m��B̭���n�w,"<Јn�7�3!�E¾��Fd�S�Zu��s���!�t��T�;4�!++"�Z`)A��r<K�Iq�����,��ʳ��{b�Y����*)�FWN{�W���2(��h�5���]���=�4��1����5*x�u��;s�W�L��"Y<z�R�����-.wpV�-*%_�������k�0�Ș3�q0�ס��l4:�.6�%�S���xڙeră��ɏ~z�p3k���Q����ȂW�@�M��	�ZV�t_g�ui!��-n�X��?G!����H;��e��+sy��v#�#^L�X%�y�ŋ���T��"�c ��PR=��F+BT:����z���uG Y�zUBv��i�"��kDo�������~�*�����q$d����2��ִ9+r�^S�	��-��=v����
Z	N����%�z˭IM6`�RQ��2Ń��-���&0l�<����玫�.�U$�k���b��v����>[��v�l�ot��[�j�y	 M�^e+,B5��+g ��5��ĕK�pTr�nTYG;7�	v�8��k�� � ��7AU�9wh~(��!"��/��[B�'l0�i���P>�D�6}/��AV�����шH���9�V^��-�j,åN�RUy����+��0��"4�dfl�fd��wh���!�����M�ͩZ-9!	/k��^���+F	M
R�C�"e�HԳ�r~�T���Z����VJ�h�{[�S��1�՞��V��I�;8�?~߄��[j�q�q=#	Kq�W�9���$k�_�Y���w��1�ʣ��K�
8{�_���`[9ZX�&�o5I��O��J�Po-2�L�OYz_���@�i:�~�^ �8��-N(��L�!�՞4L_�X؋ٮz�C^�O�>�~|��,��^P��>ȡǯR�!�77�RyA���GQr7������*ؔ4�C��:�=�@�a�5^CY~hL�,�be?I�Ȯ���1X�Ӈ�%�9��ȵ8��4�6�����9��H���t7%1�҆�!A� ��vr�Y=܀Xn�5r��j�1��5���U��߈P��
y]
ڤ� �����W����3H�[��l,�Mˑ8.܅�ı��11_O%<�ڦp��ܝ��v0C+��"�v�b����5Zw�3a�'��<47"�+F�������X�e��%FRj�3�{�!� �s����h��w�{�!�ֶ^��lzm���J���z�>��U�����(q���|�t��]�LUI�Q�۷�6�E2��@ ��~�T��B�IBiz����M1At@ŵ�ҟ���-� �d/���d�N�$�l��t�7	�`��g��n<��y�@����T�O��NC�q�O���cP�n�w�m�q\F���ֻ�������
2.H:y}Վ�p�|��J0_q~���*�c�iL�p�2^�y,��u��{)o�U�k�(�-x�ۀqM���D��*�-��oN[M
דZ��b�W��$�}}#�{�=�Eι�!#��`���B��t?�S��'����G����,���p�(Ǭ=���F��:*��0gUn[�v�F���%�4��
���F؏԰R;ܶM.�
�(�'���؁Q>����Ipu��'�=\ŀW</r_�#mCa���n�p����r2D�U,��HVoX���c��BBD�2Ay@��e��C#n=Ӧf9q��L�����!���XC��&���@]�D�W��̪ ���	�^����?>�b�'�����~Y��q���ryX��w��:ˮ����Q}�3��
�Ȕ�lT�V�0=~�J-
�s�t�ڐ����چ���(��K60k���ǁq�v�V���M��t�E+�`���㾺�긬��~	�H�^�t����oB��������:�"�
��Ks~1��}bf-�ӟ�g�{
W��!W��>RK�e�^�!0���O��/[Yt��� �Х���\��VAz��|�7��;é�k�ԇ�滸�;����~��.�zl�����سg䢂DY,1�۳<���,/P�"ws�>���)��
�����WL������~c��r;����-��2�-7�ƫ?�xlfT��O��`SmB�N���}*�n�#��4��5~z��EU{�r?!�w�3��FV��)~ �kSa��'�J x�sT=�Omf���������c���c�d�+[lY�`�b������������*��n8E4���x�B��
e�'Y����w�ƿ��w`����Gq�;�)�����c@E���Z�˞O�J[�Z�k�4�Λ=d�	�t�%���[��E��z���E�W�X��T�2b��2�,}�0G�B��0�sV������@8�o�!�)��mGs\r��m�"��n!^Ca�t�O4-��g4��CP��W��۪�Y	�)��B�ۗ���%T-��@��f��߼
cmC�A Q�[�6`i�e	�;�P	�g"౻m�q33�Y7�̂'���\���E)̇ON/dT$��mKۣ%�����C7���=J�'e��F]� �_���$h��,؇�X����V�Jwz��aʥ�u�'�}�m%{�9�jnq��~����
GM<��j�at���%��&�D,~��<&�n��Lގ�M6DIo��D"�cW@�K�C�(�()�q���tQچ��'� �C��U���^�R�&yn�@m��s"���\�]���f�~��P�+NV�ƻx+��I5�#��� �.ÁD��DZ���*Q�h
C��0mđ?����\�~I;��J�����"e)c,�