��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
���>{:nޫ��?��P���kI��n��*8��\'��u�uo,�9jJj�\�x�>SM���0���\�0���'�_�pc��j��a75N���b�[��ݟ��&�"���f��P��j
�aDa}h���n���j�BVI1vQ%�m9*��Y�͹'�u�x}�= ���@����(�9�HRg�G�B�Þ���$ףOg�]�B6�i�S�hX���Y�^��WX��O��,��v�u��j��:�6�wC`��7W]��P.O���DQ_?�����zsT1���Hl�=5�g��� 3pq��+��Y�S�ƫ��:7�U@�}��l���'���� �k�N�y�mo�w��-C�ݰ��\���#��(���Ʉu�Ub=-�������K�!ܪJqU�\C�s�to(8U2��bAl�}�^��l:�
D�5�j�T�W��W_� 	�.q)�SD����fa��-O%1a��k}�d��Q2�ŋgUK� P	�(t5ӛ~v��K�^�|����A4>�$Y�l4DV./���[E�}���Y�
��y��)�x�=�b�C^����^1H�^��� ��Wl�i�Aٱe�>_`9I[W7[?aL�NR���f�͟\��J���^8�c��Ù�c9'Q=Z�kF�����#4��3�>+����4�ёİ��#�DT<'�|��i�	�����{�����M<��޶�қ~JJ�rst�@��7�K��ʩ��� u�t���.8��*-e�`��n��	Nu�~I�\�Brd!�`}�3`�U�.H�x��N*G�v������@�a#��>��V���>����u������en�xD�O��&����ȿ��Ķ���@c�����0�s�LE���|t�〙|u�kWCE6��������R���Ip��O>�*�C�m�$��� ���y�a�"�F�)�ϑ�F�3|HF�ǵ?��V��%R�jp��	C�z �4پV�s��q� É������'�����;�b!��ΧΤ�������/#f"O��m��c�S.m�Y��\��?'g���t�d��d�d��"�������7H�+����C٤����K���{Q�#iG~�2��A��#ʲU�I��Vg
�������7�?�g�4||V �w��@)0��$䲶o��� u�8���d�Ղ�F(��慳{ ��z#5c��R�����>I�A}�9��'��?Ϥ_�
qlv��x7,STN�E�[���( z�q��nT��k�k���N6���<�H����R���Iu7�_� Z��ۚ�B��'DV�F%�`n)�^ k���^��IWK4�����;'!VBK��x�j�k����c��c �c8�½�r��d)�i������|��7�������by�|P!N����R�,ڏmO<ڝޔ�5����_<64h�S7�G������ݶ�H�EKK��<�eӷL),�����`f	 �D�6d�uD�0��J+�
�fyާ��q��\un�^N,'<w�l^�N��6	X��8�݅�.%l@}�8AT]i����:G�dbx�<���#������{�}��i�Hދ@u	к1��F�C���k�^���ԘL5�\�|�'��Kj)�A^C+�x(̧9����_����$i|�]�N��=(�k�#��q9�+
�^Cǐ �ײa>;��2X�k.�j�D�o�|�Ѯ��%�l4Y�)E�ဿ)�d��<0!��%-�(��O��4�t썃.`M�p���|H]�Ƞ�鬜�0�&�iS�c��DHca]"�qw|,%s*F,�*�<�>AA�"���/(�MaT*s{1��w-��:;_2m����]�O���	�i�2�z\e2Wcz(���T�oq�c!�6$�.m�ڶ�:�X�c���&��+�O����|�u�E.�)�91�8He%����P4��	�����鲴G� ����;�&RB�"���Dm��@8��`	@�f3�Ȏ�}_]���v�Mp� A�E�4:źh�#$p�Z6���� 1^�#`�	0/�A�ŉQ.�nZzVs�z�E�[����[�x>���N�ʵ�޼��E*�����]oW���`���
l��H(1Ho�x4¶X�?���]:���%j��,l�Ph®��U�=�p{i�1��A�t�@vq��X9^�
Pv�0B���K�r��hZK�f�6��%{^ �	^z7_���cӓ��?�uH=��1���r��)���c�dmn2��u�;�wZ�I���,٘{�1Z|"4F�͑�D�v��lzgv�y������,���$T�+�I��>�^-�iт�.;���萞+&A�~�2���q�~��F.�Q� `E�@�ً㴁r�oz,�C\�,(#(t,Mbʶ��Pǋ��>xH�u�@o�1��G����qsuY���	~�M�{!��壱3�Xg���`eL'7��.�֯2� #��D�b�N9)��iӱg��������'c)d����o�bO2ި���2~��'���R��`�ST;����V��cFW0S���J��?�7�F
�+��Z�XJ��A;@|-�L��RU���{G������gga��uagM)�!�1=ٟ�,��k�+կj|�f���؍o]⯭ڼ�b��}�v���`9B����qI�k�l�f�cȞ�'1�"dt���L���`�?#Vd�
4���R�� &^��㜱����z<L���bd�S�<=�ɦ�N��W����e��,FCH��6"t�p��/��M_�cD2�m��T�%F�Wk^����7�v?�T���D�Y,V��t\� ٲ�.?'94�E���@� ��$6�'�j���o|�� y�C댩v����M61��}e3�����S�B�A�>��E �o\�B:%�;p��n���;��NX�䦀���/���w�� D��*�u<ڡ?QvO�v�?fk
�Y�?n3�S܄���CG �3]�s����sd`�(�V�	������S^�b${Wf���I�&1��4�K���mr��^:�!�57�t�p7��wX�:ڮ�l��x��E`�._�["��ēd���lK�i!�Ц�]�:��fچ]�y�����e�։p��̼��<4N)-�&�Td;�m �p-I�R����l���d'�%�S؃1a�_xn��'�� ���K��@wK�\d'9�D�
r�e����\pEa�D��ر������D�N}�Ӓ4�*c��!b��5=���	p���X4�v�B��b��\���*k�ѠT�y����\�|�r�DX?��]�.ۭ�(�w��E���2�Q�b�nh�=���G��i/�7N����å���au��`G�W����)ї:�n������8�c�A�;�X��J'��{�+��
��d�}����#���r	(y��>Q[���D�\�38|:Z���m���4"*r�F�M���L�C����|��m�܎t����l�U������[��	ّ���ͳ
����	��t�jԞMJ�ψ���K](��͜��4Μ��'J�-����wV0�����0>�P1�zC���}`�Y��^��{)�z�}�H�w+�Z~d\��5!5�Mi�҉��W�*�@����1�Ee�v6ګʹn�uϕQ%I�Dvg��ٓScD�������Q�/������a�m�7ؔ���f�ãH�=;-�wyP	�L	׸:�o����J!��h����*���G�91����I�*l�8���H6Ă2/j�ڣ�~P-�GMݧu�Yy/�����KR�[��b�ny33�	���u��!�Y����(1^R�昆ڔ���ߗ)"�P��m6Y��bb�������2��Ce�Y�-_顷|�gn��Ov�X�{�Q���!U�_X�ى�iz/�G��΢G��m~f�$�3�f]�*�_��� �oUk�7�2NM�eݬA��C~�� �uOI7t�h��	�����^�K)1�O:��ѧ6z�k���G �E`��z�p9zw��4���kiF	�n�77��ӵ��)$���I��C���Rv/���w(' �.��Bz̶�e��{|:��D��:�<�k�s&8$���݁v��]0K�0�f�wML��s9/��@~|���A�����|Ca��d\m����%�u��*Й��ư�3WV��v1�&��a�?O�k�u�Q�_B��m��܈Z�u
xi�z橥w,3o<�R�ᢱ�x)Pe4ZG����.(4^#N��Ǜ�b�;C��Ě[��0�ǻq��[v��y�/&I�����)2�XE��i���Y ��YZ���j4Qt��Af�l�|^@.�2e���Be��J�̮j������V��VPyoǹF�(���jR��I�v�]��B��a���Q7�EV@p�/#B~�M$����g?\��ۚCi���3��9W�g��k
H��&��,Q=(�5?D����k�P�.Q�K�]k���{V�:p��`kG����IGS��(W�r �BY-��j�;��*:H:��u���vQ��4pث/������1Пy�JiB�kܻŊKO���B����Rp�e�@c��u�׉���j!�N��R���w`�V���wz�7k/^ӹ��/�`�ֻ��|����Ĳ��O��"61q:���7'i��<�Y�`����N(X(F�~ȣX%�����!���Q�'2ݾ���p*�~��#��§;zu��*�=��HTl��9���1x^�K�D�5�8�h��~߳9���f���Z���T����
�mL���X�<d|�+3$I���苛f���F�ܓ��x���e��3�z��?���� >Lo� Գ��n����\���ArN��8e�o�����F��4g�ȘuN&�L`���Q��YR�%��Z[\��|�'vJ�H��<�f�@���/��5��37�4O���
9�'����L�?�N&n@E�Hn������ 3L��ШYv�]��@��J>ήN��=�&�������2q��y��ҏ��%�g*B�Vz{�/�Ґ��Ҟ�9A�e���T�x�$P�P���{�@�.��,��k�;�P�!��m�����8b:�h���]��P=�j��)-�l����w9�l'�Cc�1����0^�C�����W cD�1W��<U�������*x�g���+{��V�u�;W�ĳ"�g6����7�R����}��m�\3�K�-���M�u�I,t~=r����ke�ΎnG�<��s ����3.��MV�9}Ȳ��m|��P�IL[�k����2aYyg%�qu����hG/q ���l�iS%:�ܯ3i*k�л$��*�a�����[v  p����I���_���W��=`9Up�禹�V	N���=�LG�O��MAQ��+ԏ��bN�JM��@A���X0'J��[��Zڠ�֚|�YQ���"~��� W67sPU�>[5�X,b��)ܾX����]�	��2�Iw�.k4���ȁE
c2�q�c���Z�L�ҕ�d"J��xɝ��v���2������D�c�����i~�$퉯�&�'��1��$��C�}�\9Ե�T'qx�a6V@�/�"�e��[���Z��X���	����л5��6��@�	���A� �^7���4ڳ%���
�;��n���fw�A�p����昅T�4�5�8���G{�e�iW���	k���6X:I�ֺ��A�5 ��܊���0�&���-$-��l�O����P��ʍ4��^��%�����9|�4$Q_��M�O��f|�	R�
���v�x��*-*�v�h�\����K�p��E��:�v�J��z1|��A9��tY�+��%R��i��B�cV���d��Z��,��m#U�}TC|�8Z�?#uu^[��T�v-_���\tS���9�Z��'�2	)�xO�|�l�ضu��!�-�{�t/��)u$��`�a��K�0�c��]�Q�gM�3��O���J]�547 �i0���<&Y��Y�:s�<�^�QG+x��N�ʰ�jg��*;���$%�y}���/V1����B��=c���/sq��(���)�a~�=���%n++�h�ǭIK�_&��{�TV��F̼3�@��н����"z��<iorHG������O��H� ���᝽��u���8�Ʃ�i��4�-���B�'��ҷ���g�Q�vFoJ�f|�����d�l�t�ev�K��6���?�H1��MU�ў���Fm�5 ����O|�U��g�QL����Y���0��9"��Yu����6��>�]Y^39��1N2����I>�`=&��avp�3��A@NӚ? �ZI�ϦFuA
��eĆ�	��S;��MN�����f�.��������U^�P���?��d4Ӟ��q�!�`ݒ��������vxvM�ϵ��u̔c�[�p��$�F���2��6R�#J(G��m�����4���c1W��dP�w=b<*�/n�c��u%Uq��u�n:�o �꛷�{U��A���*��OS���ֺB*(���P��q����+�����dĲ3�a�l'�|E��gˡ��N�����L���b�6���[����z���^.�ЍMF���{||�'���F�|���/-D5eܩ�㡒ұn�'O�S8����>HG����^@V�L�)v���V�e��̓�������	P2��B%5��m����k�����$��4Ǉ�}?F���mE�G|�H?�U�6�`�G�����[�y�\5��%�ף�O��/��Bj��E�bU�3�h[�zcŉ޲O�h(M���z��/C}h�FA��`�L��%��A���?:y����!˥��{ᇡs��`�XP7`���d��u:xH]± 4��+m�������y�^�	�;��;�p�N��r��O5%���c"����Eg��!:3�)ە�О��z�
�2%N�:��8��@�� �O���)ϕJ�nтu��³J"|X��� ����Q��q�E���ϖbg�pߝf+��GH�7'�2��)��OI���f�1�g�q�/��R��՗�b��p�	8Q�OR��c�k�&?����K��B֙p�pj�#'@:z.j���߀G|������Tk���vm�s�hU!W�3��ĊSHj��I���-�+wK��s�ly$t����
k��y�O8��/�z���}db;(��,�3tr&�ND��X��^����3��F����	<���r�f{��Ё���ƹϝ����^�\!0����)*H�" ����`g�\8�_�A�$�3f@]<�v�Èmy����3<��I_�6<���oD��!��}#Ѭ {{���6G��7��iД�Y�%�vЙ/��	BFz�RQ�BlG��� ��c���E�]���XPp:#洏G���o��#�-�{`pR3.��:��Ǵn[��\��,(y�r����Zl&��Pb�d�.f�� g��E����(C;ȃ\n6�ʔ�-��L�rՏSqچ�x{A�M��+�)�Bh7�;�=O`N�j��^=lO�Wo�4��]�ø�ɸb��~Q��o��{+����>~WQ�4/���`Hv�Q��8��8�YQ1F���	��*zYk%���DQ���ԍ���]�jH���ب�V^�����]�HD���WM�� �"Պӑ���s	p�S�������a���)�=JIӕ36�h�)�tૣA��]�U_���#��qw�#���5,�,99KWFX����a5h��v��)�A�kCF$Nݪ��Y��j*E��Բ]fX &�A4�]�jOo��N�^�<�6�l��5��d�5�Z��}���m�@�c�+Q3��	� ��L���[�A�,��V�>�jd�J.���!68��"i��"[�W�����Xl����3�dʝ�ٱ��z� X��n.�d-��C����o8�[�^0W�M%���u<!�B�e{�� �R���5��d	�1����F��I����z�Q�/��еQyo�3�	>�������NBK�B;��s��r����=�GV��B�K>D0�$5��o	�q�J�}3�Y{��[�"$�h����?o`���^T�.��f�!T�0f�O��fmCϊ����V�^��P���a'�v8�(��Gjisl�c��c�3Vɟjr���m�cwy��kt�,�d1�:?�֨)�I��3B�c�h#��v?��_�jU9�BZNQ� CvӔ`�f-[��_o�=�ۂ1l����xq;��b��"�z���0�x�h�	M�~N�.���Ck��MI��כ����=�YFX@�����x}�5�M��&�O���YZ���祚�x+ɑDʐ� �ے���� #�+��s��.Q��qh5�;�O-�W>�I�s(�Zȱ�O���^3��!$_��a%���fMa�(�u�5��q�G�nQC�'̪�Ƅ�E��D���[�3���9Szh��}��Iǁ����ZK��w��)���e	Ώ:��_����-��w���H9�4A�M<���o �cgZ9�r�����ms�,]�i�*XV�9�v����S�
C*�;J�mnG��G�[8���]��oV�z��''8�5A:����|���:8m��je��2�35%G��X��� =�ޱ׌�-�p׈�a��x��U�1�v�,�)�j2������AD���Bi�u�����H�+͆	�T���!9����Z��%ES���}M�.F�}��j'[��]=�C�u_wRE��i���N%�!z���1Y
�ES��j�s�jH]�;UKk�����g��`��Ս��%t��..#)(���V�Fn�ʌ[tz���Wz�/M�W�( ��<#��Uq8����!�E����#�|�Î�07K��d8hʳx`a.H6�Vb���ӳլ�܆̐��7�?��"��*�9��H������O@?!�RP���cU!f:��6���[���N��%t��;�lW��k�Hw͂��l&��B��
x���=����5y�qcΆn:�b�v�̼�oH=�},`�	���H(�QX~��		^@	��@:ΆͿ�di5���^2&4RƗ�s�M�yS�j��� ;�)tAm�&>�Ⱦ`\��+�������hs glΨ�!v�kI2��{���Z[� S�Ž��/���N���������R���*��� �}7`��=������(������?%��~�d�!��2C�Ư@`"��F����d*���L�7{R�]��*͈�a�S��W��h���沂fK��U�ŽG,���A��,r,!�q�R*��љ7�i0�[�'�(j9�ȟ��K�kb�X�f^�f�_/�*��@�ў0�jt3Q�C�@��b�/�Y�zɇNO�G�)sߛC �G�Lqb�@���Y�#k��V�{�Y8�:���H�f����X�I�1H*��,�k#;wQ>x3g��K&�;gI)��}�E+e��a���*Z����)�տ'_�ssj���K��������Uzg�E"Xe�6^�_�ĝ>묌��Yp+
v���9�������ٟ��/��@� �k����[�>���L��#���f��X��X��̶��G�[�l����i�?�s�KE��ǧ}"���vN��K+�O���7'0J����M,�^���Q9�]��A<]���M�*���*�`>�X+�%_��Af�%���q�)�;	�hA��:{�,�����:���+�2�y�ݤ]��]I�M�T����9�Ә^�1@�A\���ٓl�����B�����ݾв`E��R���^^�wТ3��U��j���g%�'s����.�jy�F��E��M|I��I�T�r1���ꡜ��Y
��ú	��� ����$E��u7����֊�Awŵ��WB���e�w�Ib�`��j�,����j��V#�m��#�׻8�싹�\�_��v#��3�1�dM%�*��k��ez�S>�kH?���旼%)ps��Q�7�Eþ"j�,�bDb�p��qB[�c�8_>�����: J��8�R[���w;�U4k�
����&�Y���� ��z��L�����[v���P?V3p\��f�FH�@�f,����T۾��M3����c������)���9J��P?�r�lPQuq�eq }��{)2�i�2q���S�D5B�?}XR6(�*�'�~���U��G?L������6=��飃��>�Ć�K�_�(ZES��S�#8�I���Z�^�w�*P���J��k�#����i��/�:�f�qK2�\׽�u,QK�8*�'	�f2�=:�ZiK��F��F�_��f?�!���cUI�i��؃<��J����x�tC��'�S�"�]p>�J��@tk|a$�?��G����;�}x����O'no\���\iŀ�����"Z���{���y�:$S����:�o��k01�����Cf�����H��|M�y��:ҲׄFo��Һٻ��
Xh���=a-{$ĝ-3ച*k�.�J�^YK�����%VȆh���B�F�kU�^d���~2�SxZ(�	�q�)I�b�~{�9��-�_/W�)��:n		���g�鴩��͟���xL�[gF`M8�6حj,Ƭa��	�d�tR}��M-ъEa�J(6E�!,<ݨ�N�N|�#�(���V�)MTܦ��H�|�
șTC9��� �l#��s�x��!Y��E;ۊ�"��^k�b71i�����xM2�K��$�ں8���Hg�e�ATN��
�U5���+;	Ɗ8�����h��l�)�C�ڻq�?Ոj���29B!M��6�b���O��7��g�(�\x!Kp��-�)}�0g�G@u�-������Y�޶��nI�l8���ik��; ]�]H�����s�RL�՚j��
��0X#Jb��M�C���S��7S�w\q���k$��XfEc[�f���g^<_�m�s9�� Y� x��d�
f�_�"��R��Wg�o^��!nS�*K�E��� +Fu���%�6p��9����w#�@�z����Y����ȆH0�qe)��{�E���`->4Va%�i�oDNתR\r;oj���4�a��plB}Ԥ�B��F�Ǜe���a@�X�]Ddx(�)�B�`XJ��@)��#�Jd���`��; )�&@!z=�0��cN�`��!��	@��#y�5�&W�ulG��ICi;5��#x<����V�i�k�E��S7S�L1�����GC���8�t�@7��}��);km�[�ႍ��k/�Bl)+��KX��Q4��0{��?�A��'B��4p�4_��U�������f�c^S���)D{�*������0'	HZ/��租˩��:�NĽ;ZEe�<C ��:����)~]k; ��p���dS�7|]+ێٴ���L �B]X�}@ċq�X'�]�'_rgEO��b��"oVo��]�n��勒���ք� ��S���s���H1�S ����_>�mX�\�粭��G�y����Y�3K��$��P���NP#�h��L�`�����@���(9ưl{;�i˹S[)���U���Mɫx7#æ1sD��?а�Lf���;��Z0Z���q糗�3�o��j9ا2\bN�P��JQ�}�6��@���B�o�h�.�¹�Ҷ�Hݭ^�}Fm�Y�-jL�{^{�O@80+lE��0���^�����7�@ᗐy���8p��P+�d�-�2��Jj@����L�w�Vj��11np%#O4�����HOzosb�Q)SC4��f�8.7��y+���
y������S!5v��\Pc����k��;} {�>춳��xCi�Hs ���du8�֤y_�c�����=N�]e����xc>#8X��cc�l5�wV��n$��(Gܠ�Rܕ�h��~ȳ�|��\t}�B�t��\�������"s�Vv-�����,�z���V�bB�e��KM�j>E��9R�-��!���ai4���22eO��ffs�f�y\Χ��;2�����$L�٦�+���������9̎hJ�R�Ϫ�;�ڒr����'�2��x�F�����Z�P�}��q��w~Sio�*V���3��!ޟ"º/$N�(Ϫ�C�i��L���fb|C��iB��P���x��5����o�"?��dE {��0̸^�c�V'8��M�ſ���m'��N�P�2}��ɖb�H�\^���^�~�#�0�0�֪��L���έeߐ8)p�+�O$
`V�B��+�;c�s��\��s��8��)-eZ�)*�~Jq��=X	�sǱ��uB�r�|K�V���,@����ux\H�����'�eS)�'�`��g�ɛ�g��' �N��\�ap<iJ�_[d��-�c�ӧ���{��b������,�725�*�����P�{�����ҏ���w���Pe��H�qJ��YD�Ё^X��ҧC\h��S#��_qZ�:?d/e������._��2`ͣ]\�@��2��l��?��Lm|%f��d2F���'�������at7��-)�; ����3�ٍ4����)�u�;5u'c�',�O���ָ՗��/D�H�\,#��G�-���,eܩR�\/���́��31�D�S~wo�&O#9��o7P�s�@1<�\��,��&�U��*t�x��h�E�iD�����T�F�3�^$G^m������9v �Y	E���`@�C�#e�믇�C�0{�e�)�Q�7Q�9�Of��[S��fPMx��H��?
O��d�.}fx��…�Sc���"/P�����g�׻���~�3��!#<>������s�ԥ�-f�	x�$��rp�G��h�^���mъ�������נ��Q�,��]����T��t9rқ�1d���Ǭi�~�����[`�?���/bw�y�����������Uv h��ڃcMd{暠Čˉ��uJ�W�����S�_r��5) ��	�V$�K�\��`������}�6>�!C���V��Ui�Q�NP��ο/,+�!�=��Y���%y{�.aB�ñ��5aQ)ϑ_�K�_��I7��y^&�U=(�N�PDkυj��!]@�qi�H&�P3�Q��?���nJJ��K�c=(�v-��&�Տ�ڱ<ar�j����n�����Js0���� ��������
���K��m��1�GY��ˌw�#�GQ~
2���ϐ�Z�bk_�oZ.ɷ ��;���Ne�兌����?��j [S�D�5Qi��!D.�ro��� 1>^���`��9=��*;��|��Ƞ!G�ay��1|��M9�?��
I�0�vt�����7��=�[�dH[��䆬O��{c	}o�I��#Y7-Z�����������ML�*-���%RiL�Ƞ��ϪN��#,���k舂���!��ʅ���]�#�$k��b��k�L!���pߪ�dl�|F�.�-�J9��*���'܇)�GGW��Y�b�d�����P��w�Ŕby�q�'��W�z��b��1��Jr��Q�ys��T�0��!�8??Xnl�輪|�,���]��)
��*��Etj�}RMڹ,���3��g�|rLC���ش񢩸�]��h($��(�K�����~g�	����~������^�q�{�ml��s�'�3_F�	X�C�L<���tIp�&4B�n�����c��)��uO�����*��lY)U�ɪ���+}�d�d[.W�Q�l�)��Vhj�xE���z�G^n}�y�=ϲ�M��]�M��V��Y�|vʯ� ��S��l�%w��YS�������W:c�b������=N�I\�;T7q�dB[���%/E�R��l�2��)�i}����M�v��#QĨ�GB��/(�~��<w	�A3�+��?䓝�	a�rØ�"Z���k%2D���>���%������Z@����Eg�=�p�s��Bx@A�P߅]�yTBx�(�t�_��$�JSR��W_�7�B�v��w
���wBߵ�pr�R	62������Q|-�$���I����B��<3�Qp�[�Ov�5x�&f�!Y�a�=��� �bԺ<�&i�XZ����A�0o�4R7.:`b=(e����pn��\�����4�{��^����E$���U
 �iO3�V� A��)e��^_�%���n1�3�7AeA��K��CyN��e?��I�|�+����X�Jz���`��{ݦ�R���2���G�0]�Ց,D�f�f �s+���m7g���	�H:��-$A��etn��xQ�<b�������z��7�XeI��'#�M��u ��j���m	 q�\�gՅN�q�E$���W��<������m&�+���t��r�����cE�C�iK���D:Ka�ApM�a�P� ���;�hĨmd��n��ϱ�����UE��?6y��7Am��l�1�m�D[�s.��`/��:*��L�. �=�u
[)�b|���l�b�ڝ!DE"a�[LjH��j��"����KN�g.Vp^�wj�z��_Q�\Fnܲ��]�֏DXÐ~r�
�3d��cV�	@8� ��P�jH�B����wQ�XճJM�U��w.��;q9���W�d���L�T�#��?�m�#L;�x}'�R��<�`+�:�y%rA��$���� �Uo_Ubuw��zݼ�L��h�Egx�K> 4]8A�7 q2�Rz#�8���LH�;ct4k����b���Z�c���@�3���?|�`�q���9���+�w���Z �2�zwe���c�4�SX�_ޛJM&��p�x/�`Y��h�y�/��(N�Y�	y�[�)��JWۖ~'A���I}����ZXT��-Q�)�]�t?הG��ܳ�+��`�sT7R ��@��^l�������q�آ���Z9��� ��^�A�^|Čc�Wp4]+�;!��/y�4#qg*�7�j���;G_E%g��dL�gr/>+ ���򁟺rꄽ�Y6���?�̊M��_�D�u�@XQ�����Y���CN�ow�}�U�Zi�!�<��&._?r!��V� ]�!~��)�F���i�	}�"E��R���L\�,�&�l��������L.yl�o�d�H԰�^��҃x��X��쳭��N�DS��	9�8YɅ-Q۫��h�g_\@��{��p�3C�=���	�v�M���%�e�c�qeO�}�����,EI�?\�W��R(�i��l��+*r��xjR�J����[5�;4���	�heW_D��$ԃ���c��g#wjR5'�5�.Q�b0�'LP*�P����S��(�	�hq]L�6KN�Ig`����������334CM��ި'�S��Tm~1:y�tq���G�b�Y��V+�Gùu��d���?��y��hkx$��Z���Z��UԲ�={;�ю�13@�%�ɣ���g�?%�*�k������]�������z�]��,O5C��CjV��n�.���On�1<	�>m+�׿�kF�*S��{��x���I��s,ԉ�E�r1%KDZe������w�#�zB�G8����{�(��G]�����zPr��l��w�v���q�1Rv!�$ �aE\�S�T�"Ը�+��y�E���P�1v����o?�c(�D9g!u<��?S�����Q���PwC#������;��W�1�Y�T<��s�0�Ʊ�oA_�E�фa+�~F�/Zgs�<n�w�5���d����g]��?�P���
f���i�kd>w�Rz�.����7�r��٩���x�@k@��6n� j��a�I�h'�����5b��f|�N�P�9���]�^��HF]9e� 3��G�;����Q ��ۿ�����mٯ2�'���֦�.T8��e��:%��
�w�2N�&o���5o�,�0��9q~���Za�0G�B�T��B�9V��?��Y�Ȟ�I�B=��������pY�6��G|-�TA	{1���R�a:��ni���ae�de^�:.=ӓ"�q&��Qs�运y�M�>j�"nۜ�&�_V�ɓ&
���.od����X��s΋������}w�?h��'}�r� ���M��!CgX�`��j�pE,����_6��B�@����f�����_T�cc`^�g3I��I���(%�G��n7q�qp���r�j�{s��(�^'`��= �J�Z(|�5�w�H{r����\}�6�a�P�ʗ�_߮Y���@`�ŴL�1�\.������N��f��a�}L�sz�?�b�EM�ŏ�6�,z(���_o?��P�F�'5].1,w��,���`6!���ږ�,&�ʺ�*�:3�@�pc�����5���D�!'`)?�|8��^�Z����8p&֧���Nay�1�>��ǳ����_�l!�����m���p,�Ł*n���c1�w�qG��=s��!�۞V�r�� �n%D j4^(y<�N��m
�e�_s�'�Ӧַ�C#?@ġr�C�pk�wD�l��������|���?+K���N��ɵfWMC���p�]��>EH���Z�?t��/�������E�O�G��%�q3��{N�[�'�ޱe�4��8���nxp�Jz�)]$e�e������G��:&���},���9����9�9�4��y-9!�r������^_�c�����o��35�s;z�"�����T��$�z���o�d]�,����dkK2K�}D���T��������H#�&QPA���D��E�����laU�7�5-f�d/��V$\����~�x����mG�n3��Z��J\O�U�ѳ��Bb�F�1�/*��uݟ���Uݎ�)����Ei�O[WP� "l���2}�к�����s�=�4m��Q�� �^e3���z�
�0�w�d3W�u"�� o�5`}����l֞�y�CA�G�ө���3�$��~須g���s1�
BT:$�3�S�7=�W�����Nc�ƟW;��m��4z��.�&��yF�9Gb�ϻ�g��`��4ʌw�Y��ƫ�����/��W�MH�Si�ꂖ[�=�*�,�rr.���h
��*C�a�_Z��ta����V�e�_���DXD$�`v)-��u��[� ����v{��w�ˋ%Z恅2&��D1��^\�\��-~,	����rܶ,����4J���Im��Lf�����e�pf���Md�g���8��Ճ\ї@�0sp���o�m�Ws��b����͞\�珈�aV�!)���	Ą;�̎X�b�y�%R���xm�w�ܨ�u���0�yq�X�?ŏ	%�YJ:/�=Mm�#�$�ZC�2={3n���v9)
�`���M��6E���!T
��a�[��WT�]� _����
|��)6�%�ڞd��0�_̴�(��d:Sr��EUc�HQ߅�J�e�^MWŬ��""�X������s�h^�q&G���O	F�Άd��A�1��M���F�늰��P�Sɯ�a$Ѳh5��{d���E�~b@C�磝z!�p�͇�W�������Q��*�����@��Y'��(�@�j�1���p�6���Ei�� ej4��K�5?�t4�����qo�I�K�E��\�h�\x����gC��Y�g��`�+Pr��e�V�F�v�+�O��A��1>��k_mu_��[\N���&���#�ݫ��N� 5�wH_\8�<�Ӗ�����3��U�	�r9��gW9��?�I&2Fa< ���1���u����_H������j�����}�O��W������k�2�h�)E�:��[�� s�ꅕu�J���F�8� })���i�����m��7�;�E �CO
׀���d���G�"�����ݻt����*Đ�<T���8����?W�ˎzG`K=[��n�0ڸ ;�6�9���*/��EJ)�dwVz�<��k��C�����?�3=���ڗu9z�� ��|��7_��M�ֹwD��r1�a��m~�n��H�ܚ����Ŝ0��G���[�ȃ�]|r���=ځqW!?�`��_�A�bc�j����71I%���g�)��T<�e�
Wd�?�ǯ9�߅��(���Z�u�;������Ek���ҚԆr^�fT�'q��ު������<�t�V+��گ(�n=h`1����4����X�L�V�!B��N&��	 ��ݔ�k5a��,']Nܮ��;L�!�\�ʗ'e�I��9�|y��1ß��6��K_��o[�[ �B;��K>�y^H/� ��[�<��xN��ڋ��P� B�C�̂I�4�I~"ZsR۬	W�8۞��~W>�,@�����TYx��}kO���1����G�ű��C���W4���a�'�k��ty�9kŴ��y��������@�ڿ LU���u�ۄ�V�DB-e���NjXh�6<�V�/�gѸWj��DF�Š\��$�]!J��(�7�JrL��E��E	�T�6�i�����Ѻ��I�BCe,�4�G9*W:,}�J�"�:�5�f�s<N�Hd`�ЅS4���1����������S�̯W2F�o�p۞yq�����@�Y�(�֪=�WI�tV3oft��k�;���aX��Þ�}�a�@�b/2	�=F�\Q���톪QM��*�Ȧ�2y.��63�u�K<#nn�B��n%��)�{��kK�s��G%O��,��,�w�X��P��sZk��R���� ��#���I��
��_
�,�M��@[f�ۺ�e��G�"kg�qo�� /ch:|sL�>��(���{�e�"�#�y?G�mݒ�oB2:�v��|�Y�j��=��|Ry���s��6|���Q���k�*�V��t {`��k��袙ʡ�.�P,J�K��z�N�>Io�<��3\���*�~R�)WI�AR+�9L����}��HI3����ǤpƐ �)��RS�x�#W����*����*2�	���t���O;t$j�x�R�y��	�.�\�W wq�CJ�ͧ����?G�F��i4x�">����k�����Z�ώ�i��J�H����L��4���_��!�@��8y�x�{�\`[�N�`��hu��X1�v��� ��G��PD k4+����Ur��[���4ퟷ��;i�������\��VY�u ? ��@�4T�H��v ����qi��VwU�x���i�>�t<O/ ���v�m��8�/@��=}nؾٞb�}K�EH�64e/�v��!���J�.4�_��� ����� E��x�3Y�,�V�k<��N���Ţ�{/�^D>�hT�5+�oD%H��5w��V��%��۱#�U�	�!X���X�� �	�9�2���߷�!z�}�qW >Yg7G]���n��֊���t���l$���;����9[R����~���ݝ\!%{����0��_�C>� �)�4�y�
j����������;V��\�)׌�9�	�һs����㪶�%�ȍ0.�D�����Dvd)�_��k����IY.�9pd˳'�>R)21�+������3n�+���5�!Y(k��v�2&~�\w1S�$����G����9�'oM�Ko5lF�-�j�D5H���S�t��N��u���J�a��W)q;���������.O��¶�Y.�Ւ���z�BH�O�����@��3�S.d���F9?���w�nc�\�޻����:+	�T#�L	���#�wm��NFmPmC9�x��m�5#PVu�����30�"jgw��Q�0Kc�a$\&Z*�w��W�����=����`7�k��'2���@�e�fyI�����ڕ�9�W���4$s��{a�?�i,P�3f���>���/J?ֈ���C���Z�8��Js�k�H���R�+��
7X���p�(A�y<��+�1OK.�@��M���ؚp1���n�8�5�P"q	c��ΣY5[�&i� �P#,�/oH6?�`�$x���뺯�BI�ƀ���ܡ��1]��ꪁ=�z�G�����$��F$�/�kw�⁆�Q��p(h��w�|9��`v��N�F%�h.Lӂ�hd�.JU"`4�Y
W��Ϲk�_+YwB�|�2'xU5~��I�|�L*B�*\HƼ$�ii���E֍�L���ހ�����x����]z��LI��3�������J��.�s %����X�m�Q�R�}�uZ�lC3�=�	�>����a���f�C���5�*M>HڄD��k��Ȅ�G��y��n�}�z�ƕ�P��o?�a�yd�?q�F��z��'X�����a��#����`��՚��~��������PD �'�z�L��\q[�I���[kS((@g��QfS�[9n��1�d��h5_;�!�.Ӯ�(��2u;0ݟ6�a��}\���8ҟ�2��>�U�PS?��89��Kg�{/��Kɝ1z���yU焾�>��F@��0Ob�s$[�����H�'a��Dt��C0:sQ����y��e
Oi{�1���Q<T!S�Ô}��ђ�YWА��hW��=PO��7-��2�˴���;Vc����v��Dh;Rk�O���շu�"���5����6���؊�j�)Ppcg���86�ɚ�,�m�V�dzZk'��{w�1����@q&��RUeqʽ�!J=�y�a�ύ��}�ZY�Z�/.}lj���O6��n�/T��� �FAs�[P�|������P���|7�j�`�5�.��	�PS����T�t��ڑ�G��U��"�M^�����׶Q}�S͒Q	L��U�r<V=�u�`n�DO��K�]N�R�+2�o���7�뻆D�S�Ɨ��]܁��1��O��#3�'�v�It%�k�)�g`�Dת���haC��K&���3 ����h>���(����x/y9�}&#l�b�`S�?��U�l���F�>�{a�Zf�`��iK��/ 7_JS�����_@-���=<�_�&�+ZyK6���i�nu͇�ܙRwS�2�Uzˌ�C�ǉ=���ط�IC�r0�2�����Ԃ]�� x< �mYw�|o���q����μ�{��'�N��>zk��R�ݥkkU��c��8��0G8,����9�2�޼.�倢~y3ל��3��5�4���B&m��������b���x�l��P}������R1�߰�h�c�ђ�OZ��Wc�K� �l��vr��}j�2�`�ɇ%���-�i�B(Kv��}-��>������dI:r��)徆�7�@}�O33$L����Qi�8[�l
�M�On4I"a��QRI�ؾzC��7�@���W��b�M��ށT�R5���[�b����ި�Z-�UA�ש���{S��%Jwiܭ#�Ԁ��M�e/]����x�ک2���C�jyu�ƻvv�\��J,ԣ����Hx�SU���&������]���^���ˮ��W�?�����3V?�B�
0�]����E�_�!Rq�1�`�L�I���I��vmwQ����T�����y�$׾��B0�K2ua/��?��su֌�>g���dZq�C��avV�.�g	�p���2���%a�m�EU�O#XVj�+��/(�0��"B��}y�V1���S�fnᲢ�@�f��kC����ٴ?6E��Oć3^p=M�{/�>W��)����-{�Ճ `l��8��ب6���2�K�5�5��[���F����,t��0�,������\@ъUX#��7�^@[33#�R�7cS�n��Pޒ���}������Yl�N%T�vp�ͥ��Ho�_?!��.���Q^��Ė������Z|k��Ħ�\6g�:��m� ���Z��*�2���O|.B`3�.ll���kٰ��D'�flmٹ��V�P�_L�89�!u�~���p$4%jf�]�rp����輦�{�Xѡ�0	�gfQQn姀��u�J��1��f2��	�<pg"EvB�d�Xi���i�]�x�0P �֘aɔ]V!E�Z�w%�'s|t��e��p��x<U��&���*"�p���!nZ�����)�rg���7���bH4j�JA`�]���+��-<�ہ&�Z����m�ܙ���R#j4�u�&kI\���ǳ��0���"7.Y���.��EK^�\P"@�c�8��o+c�̽�!��@�b�mβU��/"R]�L>�� �Uۄ���왺^O�Q��a{T\'#��H�s���!I�v�@�����,��B���& �Z
R���2�F]��S� �)�Y3�nc*�'
�,���u`�^#���Z,4�/������r�M`�UPٺ�W��t�{���%*����-Z���9���_��9�5OȐ*ƑJ�7��� ��(i���f�$��Sa�3�(+����Ҥ���osl���fn�M��B��=���蠃}+�B���lTc��P��`ʁ\�l}	|,�h+mf ��;��N]�{2��+7@>�}�ϊ��B�雡�.y�q�h�O:ǭ'�jMiBal�%�uH]��Jp�evҖ��h-�7��N�L �G(�Zk�Y�􊻡����X�f=���d����e��w�?�_Y𷨞˅� ������]^� }n���H�J�/�h7	72#j+&T$�?J`�F��\iV