��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
q1��S����5�~K� ���ˆ�AM��/S
�'�����ੈ �<Z�{o[��9���] 3�3�ABE[ԑrH�]b��/p�����LJf�`��A�t#����?�@L��#d���*ӣ;�ʹE��������u��ʚ�:�t��z����}B�gNC<��D[U���"~�^�{��&�#DR*����ff)�rވ :Fm[xa�,��#G�`_-�o�K�F��K�o�&6��?fp� ���ܟ��	�p.?�Ygg����NYd�h��Ktܪ�Q�K�R���rﻔ��MHM��΍�h�r��q�?��6� �-�'�β�YƓ%�_��М�NhčS1c<�a3�6�)�k�
&�G���z���sa�1�o���3F��,3r�ʳ����"�[Cq̼��P�J0�pNֽt`�9`g�:�g[_�83t'�?�~�e97W�s���Pj���]�v��>Z�=^[oa���o�-'���$Hr���Y��o�amثd�
�#�Ɛ5�ܻ�G�S��r�Z�����h� Q[u&�^[��$�)N/c�6ӫEP�p�}�'G�G��6'�qnZ���$����A�Z�< j��m�����vϸo��k��3g�7F�g�/�>��k�9ɼY��#__iĘ"P��e)0�����J�����x�!iԃB��+�,m��PJ�!��C����ު��;Y���7<��3��a M�rw(���r�\ֶ�g����S��g��H��͡�q#U�l���Jm?ͅ�3 ����rqd\�����KnmU �-}�&�_�Q*�Up��&�����W��A�!g�d��!�*�kk���?2���rZ��gRS�>v�>r��]`�����SG̶��R�9�鷹jhQWlN��Y�"�����MMFjJ2[r1${��4� ���%㩍Q?��34K����B��I��p��ޖKbl�N�M�N�7cDVw�wK�k;�=����l?&��؍�V�$��6`qe�h1Ѵ
��$0M"�!��[�}Ƃn�R�η�ut�O��7��2��a=�mXk'X6g5-���N��4�c0�v��g�����O��j�!^���[�1V���MM_��M�/q@�-eU� ���nK���dJ���a�(N��<l�����A�~�����?n�)�x��L"�o�H�	��-�F6�G���'��$���lЇ�j�[�O㹋p\�4�� Qѿg��B�Kh�z�Ī0�@�_V\���Z�TKB�F��~�y'3������Y��ܳ�D�����2�<&�M��:�ߜ,I���K4���`�⋚?xX��\���ʉ�[�inE5��8�
'��dETհi}��aձd���a�b�܎�8���4�Dd��ˁ~*� OzKU��dl%e��ͲtXPȄ:�V��:.��Xa�}��a�g~�rܸ�+`��M��h[V'l"ɠ���G�lK�����ݚ��M�s��v ��-�C�o6ZD<z����1�Y8ެ�������u˞�u�U�Kgې�]�����
Y�mH�*��؆���M@E�Y,&x�=�l72���J���їX�+^6kû��w�Y}�τ�#��pEg�%ѥQ��>�޾����kIu�4����y�`�4Kr܌�'�to��a�gU�@i�oD��ٱ�G�G��2�ֺ��"�?&���&{)?�����L���C��y_@j�	���Ƈ�ߐ�]���<��I!T��;s���Q��F�,ɯjQϨ
(��i3�4��n1���ڧ���K�Jz���-� ��fIzg��b�fV�L�2��Y�X QRo;�s@����S��e~���z'x��_Ok�Scil�%���aEڴΑ`��j g��ܒQt�bW�g9�{�d�����'<��B���<6b�`���ﻏa	�jc��st���[�:����BI�I �:q��.�墽�lyKR�r[&+����!�?����@���ia�j?<)�	�����+�4r���@�����ahI��-
�s�����k��Q$K�v��[�c�<��Q��(Q�M�G*�#E�s����&�[���s���*���y����Z{�h��=�S�@�չմ�o�l>ZLj{{JP�n/z���A���я���F�Z�セ�t�jO��6S�e_����QZ�#��m�����w�F�l��0y�-Q�������=�ϤV}(�_���t�V��is� �I��l	[+���B�u2��淋H �8jF�ha.�I=�&�������ъ@��$5���jl!"U��tmQˮN��Ȃ�������a�tc�m��e#T��xQ:l߷}YƌI��x=����z��t��Ľ_ȐY�$�P/�q���]����F��D?E�-׳b���I'*�w	yxHl����۷�;�����O��k��r�5ϼ��> ��-�S�I�����w�4��/��g�;F�7�!�p�X� ����0��%�L;�f~r�I��'%U�6!�q���s�-�ϻ��X��r�%�N����xVob�:��,J��������d�d��S�+�.��� ��=��"M���Rp�OW�;rY�X��KI�,�̤]J@10u�������^�H-�7��m�
wI~�3�̡��D��B�9��*S�\X�Z�8	XX'���BF�C@������;���m����V�FO
���m�q3m������&)-,� kd��!9~fa���#@P>�KkJ���u?�D����$kr���GB�k�6�2S���ʯ�'�l�^�d��f���-}C���`y�����l��)b�ϖ�֘Q�k"j���� '#A�6�A��S��9{nu�IOA�
�\��}������,8�k,�g6<�LH�Y#2��/�����&Vv{��U�N��=c|9�p*^?V����
��}��d/�ړ�����f`�����x�|k��I�B�s�6���c�%�#�%hRy.�U��nr�JF�k�Iug1N��sߴЧ�N���N�/HטIv������]�I�	��tS��0h�E��Zn��}]�����$��\�M�{8R�^�l�����nB7��;��Kcm��r�J��|
#Y��B׸��0G����� 
T{ш�x΅�*gd��^X�����|���`v���D06r���P\�`R�L���Y�p��NS݋�1��Ʒ�?��Kr��{�R��t��؅jѱ�b"�/� �Ǿ�h����O�"0��FPH+��lz�'3���Q���p�?w��Ra�Fإ���#�y���\���.y�t�
 
Al��=���HFQ��9ڣg��3��KQ���sW:�[���_T��^;��;Y5wɩ��]�IHDX3��"|��rSev�X��8�[�����]��:v���k�P�1dz��;��}gù��P��s�?�`�O� �t���E��5&�UocD}�k3��D$OE�O�oLȶ|H��S뭗�7W�D�W��0��y��@m&�c!���f�˔���@9(��N�H�
]d�s����)��㈫)>�+8\�6��-�XGD�+(Q�{b���Sя��#tH��<����
(2�;��?_UD�}�^df�Uz(��$=+�C�/>�B�2 c50��g���GQQ�����<����p!���;&�=
	H8=�n`s�� @"v*g�4�H�Ȝ 	Y��2�]�Qn��1P�~/�w2ˍm�43�_�������64Z|$]3ӄV���V)���ɒP�<=�ߊ�n]39��GFp'�d����L�':����:QY��*;���[v&��_\�/ -R���88̳�v�܁�n�~�����G���W���x�\}y�� B`�(C��$R��ό� ���������A�䱧;7���Q�B������:7u'5@^�� O���w�b�����]��	~ԪB�Z�4��SA�S��l:3��Ic��D��t�����J�鹱ݧ&��щ�D
7Huw�:����
���:&F����r��2��P�
���������0�݄Rn6 ~���;l�!/�@ �>�;�<����}��f�a^q�A���� V��L��x�K=�fb��bogɋ���9(՛�;Z�����mά��&Т�j�ō�6���h�����"�n(g�9@�:��e�Ɠ�V�<v;�9���:�g��6a����H%d�,�6i%L%��_��@��z4� ���J�0<�P���=��;��T�*��d�3��t<D������I��2��գU���o�m�ݸ����	%�N��Y����Py�839eR'�0;p+�Xi:z*�w&H�����	k�ֵ�Ҏm�J��q�5��{��ck ��3�t�������@>�*8�-�V�C��yS�Mo���~)\
�X$�d���5䎻�E6O�gR��ݧߓx�dS~�[t���4��k����=SZÉ&��f�`�7�:�.������S42ig��
���n7�(Ӱ~��w͋H�8G�y�u�عY�� ��d�#͌0�1:icyA:��3u�;��@> wD랩�ь
��v~'��
�~���d_�۽}�����7p!��-����oH����?������4�R?	�A�^���n��~�b�`�r'�iD$�|7�@f��!i�,�YFwP��pe��>�Y����vd��w��	�H�L�>�g�D�gН[$�h5|��(%/,a����D v����i&�2���7�m3��6�_�:L��֡�"��(��XD�Lx�_���y�]9�Զ;t���.��Հ��@���j���X#�=dJ�#xֲ#^<���h8T�I)����O���5Q�A���]�?������A�N���l�@�]H�Y����n}��b�}|�q�`�Z8 k7UM�ͩ�*c$�^�Uq�P�zf)!�݇�颃-��ml�q?��z"a��F��&����*W���#�BAЕ�L�W���e8_��a$�0T���9��&x&�g�x���3 eO�����z�iq�+#r��`۱V��S��곹T�
Pd
�F��9�V5G�L8EAgZ��ҹ��Q<}��Gγ��r�<NN�v�I4�@A!9$��ɿ^���9=���=!D�����ih9��fx���(/aٱ��od�H} ��0�U �x[�-��9����+T��`8�gC������DFJ}�M�>�SND�~��:���G����w���	���㋿��[�&i�mF[%�����R4`�:�;���R0d�Ů<�yExކ��49x�K�y�0Xt% 4fQ]�ܟy�J��½k�xA��6����`7�y	�u���J����k�̝��hdc8&�0�|����1�X�J-�Sh���@I�S?3+���Pώ[�����M���	_�k� Ï�]�	�O��If����ì�,?Zi�*���T�JmZ�YqI��}�֒%�/EhF�+� ���h�z.���5�E@z��m�-�x�WU��R��`��襈�mY0$��� �m������p�5��zo�s��>��;����y�Z�(_���y..噏�396VV����@Q�w��p��H�+:����^�겶�.�g�˴��+ϒ��^��^7�5����vL͔T(r
�0��d:������9�e�JA���{8s�
�/U�f�cP����YHb�d\V�[ݣ�hi��7��̡��Ug�~�'�}��i�͂
>�s��	�ش��:������:����\}\�0E���sl�ϵW��uh���+��?f��u�<�ce�(p�`��{5�B�48cl����iX�Y�Կ��������+#�P-�t6Ҙшo�u��n3��j��^�������4� ����I�X� �ʡ�R�I�g�������+-�=(7�0%�PK�2 �����a�����~�����T�����ԧP�j{��!���ѳ[����L �|gF�:!!�o��1 �,� @�>��)�ɀؑ�uS�lЀn��;�b�p��]�/ �r+�#��O6���<���������/v?�MܤwвE�ro�g��rn����{٬����E�K&o&��\��e��Y�z���n�L�l� ���D�$����3 ��Ƀ|."W�]
�����K�e��M�h<�vA ���C��/ UI&����c5%.��v.��078/�fru��YH�ޙ��	�NR����^�/�$f~i7�����6��O���z�O��Ꮭ���x�@�)� ��eϱ������G����-�'],M�JvA�d�p ǘ�[��͹��'�i3Ʒ�l�70w���V;���
�a��e�兽�H,o�i��t�`|��D�@x��e�i���_h��s0q�"©�oD�̮�u�;�I�j��
K&G�g�Ƙ�Ow��rW[�C)�cq�����o��V�h�g��~pǬ\�QD;�冽n��U����As3�(����X�@#�;7]�sy�\�`��Bb}�[��@��j ���re�ͱD";�Nz�����U$,�>�<��fE�l�4`25�Ћ��A좩�ʽlHZ��n����!��P�0k���D��+�}V�#�*��1�7!�:}�C)�t>n(~�\5���G�M�~󵭂"'�ѧ�e�pg����4a�_���w;�0JK����Pޓ}���AX���$�dH>1���V@�m�]��m2�mP�5��<Hqt-~ԛ�8%�Fŷ�N*zǝ�ţa��n����9�i.r�QI�N0߹S���X�ـ���:4�|X.�3?�7e��
&�^�T�OpCR�Vi��q��E�u��PJ�",(5��}��٩���PL����-%<��L���*f�Gc��%?�2� ���a�=��va��k���Gl9�0�WH�+�c�MjL�'D<􋈝�fr�VRZ���d~Mt�b�T�'��1��{�or@Hqy����c�C�s��fz�[�z��j�P�=�\S���>���h.9��N�ߚ[׾�Єg�{s��ָJE�L.��9r�Ԏ�v�jZ}��A!�!�&I�7�W���b��6{eMoO�P>�̵���z).`�!��`{)^����*n,�R�/J��u���ZE'�C��uU�#5���х�ٳ`f�k���@��D�x�q|�z��R�z����d���Չ�Ec�i2�Z���D6��Q6��/=N��͇��/3��a4�OZ������&��ud_u�iǧJx����^������VA�h)���ƑDL���X��&&�-���/�v���Y���v��`���"���]�oX���^�@��L # ��v�����-�t|uK�ɜ�jLz#�_;�c�q�k�	��2�e.L7���,��Cո��:��X߽�Hc���|(յ]�+T � )�K{�G(7���[�)�O\;4W�:Q�޷��[״�{�ՙ��ȯ	��/��W/H��[� �U����W��Z|��}���U#";� �4�r*��d��̆X��Z#��G�؏^�I� �I6Ϗՠ�$6�״���NbNR�>Tn�f\���-��D$���{/t�����FE����,�3�"?� ���!�)��O~qm�5��z�n�@f�!����u*��f��\�{1���Gk�A��0�S�իB�W�7�վ�"ˋ搌��g��&�#�+1P�[���GuE��R��WDP�k�Z������mm�ƺ �^D�r���9�H�]�0��c��a|]�B �1��xXs����k��Xa�;jO"����P׍�u�8�7��^5r�w�-|8e?����I�fҥ+d��.�U���ʤ��/�Ҫ5F��D́��PjA6ʊ�X4k��7#��B\��0�x<�q�oP%FKn���2�%�HԖ��1a�)���2݂]`;��`�L,��;~#~��j�����R"K��<�f�7��K�7����"]�A ����n��m�9'�����wѱ%�k`DWY��@�h'��$�kp��ŋ�)w��-�T=)ͽ��#F��Nb�<�����F11��ˡ>�kiA��\D�e^'�z4�����[<�4�&a���2��v���h8�|����T#z�v�բ��D�тܼ��j��^7t=$�z���̱��~`�Art�/����o�m�d�xWp�t]��J&%�}!�
,ukh�Và���Dї���#��!9c�&ə���x9ܼ�y�����|L��'�����u�߽��N6m޸����7�J��ʠ���``������ޤ�\��"�Q�o:H8���N:�Ƙx�R�JS���r�Z�,��|k�7�>�l���T�̋?4�����E�gEPg)Սl+ڠ_&��i�i�|���#�/Yv�^y�1*�?�������n2?;E���w�o�	����uQ��wi��<���6�~���b��AIĞl���)�g@�+]|d�:���V�NSizL�p�)a ���43	����\��=&�x|�����c�T�wU�g�r�^̖��K����R眼��������*J�  7m�Yg�\(���iu���j������}�~�Z��1�G�ͣ�}��}�.��bhf���0��f�0��*���"�ďw����[�:ݛM���6T���Sf]]��ay��� �ݫ��d��Ջ�'�=\I9��|��3��h���!����B��� ��Fѓ-�%�ڬ3�l�ڤ���X$#8;Z�����v����O�Xl�BP��x&m�
w�k%�C�&�2<�9��*}�*��oΛ·��́*��V^�q���f{�>��ܝmc��_7Ѩ�a�%I)�&����C����$7R^���;����5iΕ��4�GbC�?�@�A�<�;��G+�z��%F^������!�����O�]� g)��X� �m�7��Kw��"�#9��T��}� �T[��П)M����3�6sܩ@i������J.T>n_���c�����W��3��>_1��ٝԡ�re����*���-l�[	[��m��[Mu�=ghf�k9*a|��˄�(��&��ݫ|���TI*&�}f�+<;Vk_�%��SJgJ j�<���9�����p��Z���D^�a����F�2����*Q}������+�o�Ӛs�c�&.�0���%��Ap~Ut���#��֭��y�J�����BewSm8��_Nnj�6N��:��1"\bR75� nS�.a��ri��]C}e�@o��v#�$�8�Q?�$�H���%P�ֽ����*�:�)��b�&
v� ��=]��E+Ҥ �	U�FJ�D�x`�����h�_���,i#��8�ZS��q,�غ�\3Kf�q}5�k˝��n ��OkI8��}���Jb6E��9Z�c.���3��S�!�mes��u�l8���p�!UŃ���>��}r�^��T:Z�I$=�@H���ZaX�f]�&�a���r�6��L#d@�=r*�ſh�xj������	�e9Dc��y�`�F�'��M��UV� ��E�	��<K_�	�+.�r	,AOGJ�վ"#�ͅ�@��R�S
�0�w>����5�;�#��	"5c) ���,-jee��R�d���91����}ܑ�CK\}�f��wԐm��zO��g���.c�;�'p�t|�1h�!��������z�qd�Z�b�������}�/N�Q�������+�dwq�M��`����^@믴���$���������,�Sڞ�\E7��Yo�u�"��a:��Y"1+���Q�U�1ĐH6k���F���{��8A2�u`p��x&��bm�E�=v����	����o�$#N[��gE��Vr
s�^dE���U�}8�?69����u�*��):�C�-�)�)ϳEi<�����b�A�H��+m��r�s�/ȉ�GF!J�f�=��I���O	�J4�s���?��KKp��V����g�j)���?�4V�������&@�vv��������Wu��+`ԠL�����#a�7Д�@F_���uw�5附�0gy3�(iI�?��%b����wm��r�f7}�A��/.�]�<��A��d�����-���^"�@�6�1��N?�
~�q���'z�}㌿B��S�N��o�� i�	A��]W@S�POwuo��s����y�{f0��F��%���( )7�b+W%_�l	��o
~6�A�� �'�'�d����6)t{ �s�I�8����^�l5k���=��>u�/�D��뻢?�a_��b��������Ek2y+���� y�>V2��G����gZ���1��`�*ڻ�߂;I~y�tO�����L���MKd���
���1}H�̰PƠ�l�N�p�w��[}��ܮ� +6.0�A�I��yELT�o���5K�1nE� H: {e�cp$|��9_���<|��^���\3�i�j��y�&x�3�/��D��ٸi�F�4^vpu����x�׋I�����pQ��[��C��ӯ��M����>��	��4)[�o��Ų�����qCS��	�K
�_6"���������?ǓƩ�5VJ�F�J�ƙE)�Հ_���y'��56`gL+�Rs�%��{[֖u��u����mz�77����Ϧr��B���d���3rє%��O�A����T_^)Wc9Yތ�*-�k�pe����ʀ��5A$�~��i8��10��Wڱ��T��_����Zm����H5���՞^^[&>)�b+�,��[al��6�9��_0��`�H)$n|g\�,�����k�\����1ݿ{�b�G9��,��Q�o���k�C�zK�싏m�+��;�MM�3��@[���W�ͅtى���_N�s�ɣ]>��r��QШ�D�8mߊ1�?>��(4��֦�f�0[+ȍ-�(J����}��_+����p|*#L�X���8\���.+�Z9����{�".H@�/8�w�[�g]���9�RP�NEϡ�0q��>����ً"�9-�o�gz�K�a�m�&���<އR]O ��*�U��c�����=دIJ"n�Pֺ��P�t�b���ZP)�'6����
	{�aR}Rz��a��CM�dc+~+����TG��������Ǻ`�r���_�j�1"�:%�<!�i� ~L�Q"���&��9T�D��Nh�F}0�g�P���X�{.?1N������.�ʸu�h��	䣲��ʧ_�e~��>Y6)kN0ܔr����k�r��;��P�׶0�H㞐�&-�57s��胉D�4wp��-+p�q����ܤ�K]�F�32A�x�89�E彃�!K�#v�� x�+�T	�&���̌[�5$"��,�A!e0K�z[x�4�v2B*��550�5�=�Sn��&�^�Ũ!\���5�E��]DY�Yt'���G�_?J���#<S�/&|�H☶\�['��-�Z�qĸ~����&򳚍d� ����*���w��i��v9qC�n �~�S��D�=��Z�n�ã�+�^�`��R漦�ScA����m��d�zd���H5b�0�C=�JㆎC1�n�ܐ���"la�ب�� f��tO������%Ga%������El�\�U�?����fs,VF5\�P�k��9�N �ͱb3�/��O�/�IM��3W| �l�X���,��A�g�,R�f4�\g[�cx$�z=�����h}�Aȸ�M�kۭ�璘}-܇T�Y�j<{��bsi����j�%����(^���X�c�t	�H���W2y�(<��ĺa��Mͮn�n_���!��(:��r���פ�~�Y�,�����ݓJ'�<t�d_�� ���������]��T�+�5�^��Ү���mT!ŜQ�����W�hF�=%uj��Z�=��Ϯt!D?xْ�u��V�է3ذUZtd�R�՞r|I�ԉ���m�d#m^z������~b��K�Bh T1���5b�qD5�!D�d�A&��4;d��s	�"�e���}�+����̳qiU�/!6��<�$��Z?#h���z��OG���z���gW�g�~W�з�o15�5�F�����l�?n5in�z��K�U�0�FK��f�~�d!22W.m����T5j]�wT���t)��hw����pr�PQ`F@%�Z��%Ǩ��EaF����6�m
��h��)ٺ����4�v�����E�s�a����q��o
.���0B�������u1D�t*p�x����t�u �'��G����I��?j=��޼�X\*#d�~��$yKOp��W��������¨K�	�_B��T'՘��G���܆߃*50W�T�_C��O?��A�#�N�S��k�@�
-�%@��n�M�NI����Mg�T-+���p���4��Fq���n�Ϊt��z�Ϸ�����l>�\�a$�%��f���o%��렊�{�w���?�����*x,�K�A��n��4l�)c3���������o�|gW�]�#y��2����		��)H*�/ � <��8�"��ԛ�/�.N�'^Pr�?�O�b��5򁚌P�>���]�����4�K,��ܨ��Ձ�+�M�}=�8\�w�=F�,��zi�$t�1f^��!��M1q_����t`����G��+��&�Ń0��?Ӝ�Svº�W��XE-}���-�D��`���h�;=:^���H��p�ӅY����=Z�Bb#ހ��_�h)=I�T�N���b����yh�w�g��J�'��9��`�*h����]-=#S6As0��E�ftd�s��e1�i`#M��-���4�7��	��5�D�IiXa?�����c�`D����zPB�!f	Л[X8D��ʯ5�<�3�يjG������%|�����9����k����D�\��x�ʵ���@�Fq��v��Y�B�V�,��1$��Y	�h���.�u�fb�_3���6��W�4C�!ꉡ��!��,�0� �*W�~���XO�.v�%��ٷ|�ܫ,��J��lVC9�3/���m��"�'�v>&�Ȟ����vK.�]s�0�f��)n,ɪ#GW�>����Ն��I��V?œ��L�>��;��K�yX�Ppɹ������#91�#F�,�N�`�L�����}Fc����RE��-J��������>*���!�5Ѻ�������l'.����6���O0[ܮ9�$C�FG�[�D>qF!֌���wh�ԧ`�ē��3K8�U�5��ヨ�A��.��$�?����f
�_�.����=�d�be������i�&�B^$�3�z}�0��O�`�>'�OL�Nɜl�>/��A �joX��,T[�$�9�����V�t��(�i����(QJ�f�]�~��s�Al�?���	~J�����K��~{-��`N.�	��o�����[�j��r�{�}[��\������+myB����Z��������*���c�&�z�K�(�������n�A���gK�1 ��9�n��M�I �������E�V��ܾ�x���`��vh⿭���f/�X�,Xf�v� F�B��]}�\��}�C�8��~�"�Q:�	���g~rr���1(�+Kz����x�Z�� ˿*�wV�R�D�Q���Y��{���$��~\��I~T�jƾ�,�/�Έݏ��H��G&�b��a�:���)o]t��`W`��kG�P���7�������R���eqq�E���+Գ�R��\�e��.ɖh*xӀ���, �/7�˨��cQݓم��IFWhç~�#Ҭ��v�^@(����́�BR����t�S1 �\ӆ}P}����֘,Q��#_��O�� ��R�H���c�@����n�oE7�6 m�f}�0Pa����k�мR���L���\L/�"#J�����0�
�d[��s�Tuf+�A�w�?���S�B�4�y�7%�z�U����M��9��3˰�ҧg3Uc�>�5��Ï����a�(��1=����A �{���Ƞ|��л�g&������ﾋO�J)�Z�ﺺ�[��-��HAn�xm�����Zp�E��/�yc��kO�i���t����tf�0���|�큡���y��+t�&�E�I�[h�LY�'?�&�6���"��8}~�s�� �*�䷦v޲A]������7�e�ˏ�/�0�e^F��G�E�b�����[����g R�WEQބz?�c����ޕ?�G�$oCZe٫�Y����wTq��	T@|��'3I�����DŐ�|��_���y���&�	%wķ��j���r��a��]p�q#�ɿeD���(�0�Ge��3:�R�tտ���:��N(�t�M�iSYFH�}�O�f�	�/�Es��:~	Z�Ts �ny���v�e��m��&��7�qG�y��M
���ϐ>�� #��My�Xƒ��8q<�qɑ���K�]���t��cl�s��]��GH��^�q*QL�u��}Y�ѧ
�I�}iB�����=l�(��kw)0����Q���Й�u��qZ��$WO�7_6>ض޿u�X`��&�����fW�5+���&�N^y@^i��g-0����&��M����tF���?o�ϖ��@~�?2$�%jϗ��qP,�ޮH��=�3wwpd��H�_�a��t��B;�F��e���l��Ù�J���s1��/v�xnJ�´��*�����\�� �ms��Hg��J�me�B��0���Q־��ː�Ѵ?WYߕj��P�7�H�&�x��M�}��-?�}M4R��;�V���n�ă�ιA=�x5A'��,D���'��a�X�1�X�h�������a�zK�y�ol����OtOg�t��ѡ`��	�V2fAI�*�F"5�3N��Uia09���p�-��Q�|Y	��=�X\�:$ݓW�$XRh��Ӡ��`�y�QW��6B��u�N��\)�ui$�q������R� (�R�����bL�� �2��.C:�.�#��|�Wy����JJ]K��eUy5�^�(��ĥ��H�7`fipD�>j� ;��Jԙ)��2�y�8Ȑ⯓�+|t�_���J�P�>F'�F����v����Wk5f�"�ܗA<��G��Ș1ݼ�}h*�hR(X�~;ly4t��?(Ƅe������\�VX2U�!�9�D�k좏s c|�%���Oqqp~�v�R���sL�@����ly8¦Ih@����ȩZ�;�d��u7��Tv{�(�xrM�V�<x
@���Lڝ_Rm�9��8��_�7�(��p�*ܗ�)un�6�� ����W6:@�>f���ѝn��,~d%p'����
fA�m��&f��9��c�P�tw�_�J�C�~�ڮ������0� [�:�ci��F� �ҿ�U�� �UD�`��������z���$��L�X���lõ�����@��&/��0�Big�~����v���u����n�0�O�a����(R(�mEǡԤU�L1�`ۘ��|ND�5S&�m�TR=�<��$���8cʍGu]غ\wG��ft5XN��Yb��0W�R�2C���1r�>�'�,f����Os�F�5z�(�d��+�N_8'��<_�'{�Q���k����0��;���(˂ !�\z�nOHZ�z��#N���&��oXoNk��V�~�JM�
i��)'�������8T�lm7�Yw�A��~f2�	>�XM$�Aw�
���q��7|%�^tj��^���M��C��3�p���Lmϵ���6U+����9�ۍ����t;�O�1#�r2��ܙ�b���L�I�XY��u�Ւ:��?ŋ��p�_/,Nz�P8.v��ʱ��=�c\���\p=U8�>���
w��>fB��:�an���F8ub=H������\��-+��n�d�&��O�#������㒿ؤ�겤(������;�Ag8��E�_$;���>S�_������q9q�U[W��z;�;��"jt�R�AS#���%�比k>���G�m !��T�J����-������(�9h�?{�3�U��[�بV����U������C���{3��m������]��c�Y/B(#+�Uxg��Ӆ}q��p(V��ʴI�Iރ�Ќ粲��KJ��x�Ӳ\����iC�TD;�ߧ>�)����+����JvD ��	�7��7-� ���䨜,zG��������T���M�t@�P��Nf`�]���z��D���i�P���ۚ^�vyX�;`4z&�Wp��mE��ځ�]�����9r"��3��B�2-����C��)6b�B�2�P���YM	�\v�;&��g@<����S,n�ˏ�c�#ڄ}5�3�=��`{����9*�5�;����ᳶ���-���X½����z��{�q9��� �h#�LX��M.����2�<��1�PWQ�q�d��������r\�<�i���`�����o��'��д7/���Ƌ��\h@?����xkk���ܜ�f�.}P�z��?�V�"�g�,� �B5��#�e���r,-ϩ�S;)�������m�+��x��8Z
,�� [��e��:yxX=6H�'���WU6��P���w�m��8����S�21�$~�y/��w��o,�ʁ
X�@|�ǜ����).���) W4���Zr�A�gW@p��Cx�BG�������U��d���0q�6��N��̒W�߃'���^8%ـ�JIҋn!��s�ށ���q��.E�)�Z���
Ss������q��#����T��O�7�R(m^L�Oc��������gB��	�Pf��]~��|��2�e��0�Y�N��宵�zH���"k�D��5�j��o��Lf�"�" �m8��H?p_e��w�M�G��C�dV��s�JMJ�Ul�N�@��Y�HS�$���;0y�;#�R��Z���t�|���r���d���2-p������i��@���#%3L���'O�� ��xC�+�9�>���3D�3�6�#�X�KC��P�F���hͣ���!�+��9Ȇ���䠮ew�H����3|D�t�pi�J�C�n~�"DP���*S��z��1�ŤZB��2!�)�:C?/�'ω�y� �ܫ��A�(8<��3Yΰ
�Bi���A���>ФQ�$M�Z::th8fԫ*�Q7^�Acu�m��ݽ�=S,Bq��T�Ĥb6�a�\�Ԩ0�,��2f���>�8 ���2(�%m�i��%�^q�b�@��d�"�1Db��+�H�^\�N�_D
�%� �iO:�}T��nK��,ثw���v��Ĭ1h���B� ;G��,"�>�8�<˓�J����'\W����&6j��H�-^}���!��vClv?+R�׵���_�z���y�r̵���7ҫ�گ��d4��R��&�ߤ�ZR���A�4�QH�UʢY�:�I+�w�j����L��]��Z>Uw0�p�]�L�=߃�l��6�m� O�H����ydZhaQ6v��n��@��H
�JW�<k;w�_����^�)�Sk "�N�Z�w�EFΰ�9���ڳ�͒�diϾ�H!q�Q)��A:=��R�����DR��\��Sf��	 ��V?^�p3d�-Ըt��c��7�M#�G
�-TWb���:��������m�Gb[V�zFst��M���oZ�w,�3���8;?jlX}%@��8��Y���uQ5��_N���;&�b^Y$v���݇�$̰,�d����� �Q#jM	6�!l��{�z�6I@�}�V]R��&��_�Ô:���[�ȏ�hg����NP2�G����ٓ:!���L�`%��b��Cm����3'�\W`��"F�cjc�
Ci���ֱ�4�������94nV]��Q�g^��:=A��\=wM�d���څ�tLu�b��{{�r�nC���Z�c�O�
����,>	���z󏪦�#˂2r��%�C���'$z�+0�~��_[m$�w���k~����T+����O0}���cO2�H���f]ɫ*�vmT_�1�i�iL��gȟ�Uh�$Ȼq�SG�̅�jrNE��¦j������vt.>t�0���İlEI]w���{�U}	�İ�B�JN�ę�rN���ŗMyK�I��I�Qg��4K �1rB��E%P��ߝ��a$,�W����q��h<�$�z�@���V�i�-ױ-�[��&c���^M��(u�+;�|��=ڢ��w&wiA)�a�q�
�*"���bo�v?�k��j܃���+͈�+��Ji�NM�c�*�R7V5.�+�5��M'ծ��ҿpЫ=*��}��0s����N�/� M��,,L�	YZ( ���w��� v?��I[AQ�1�@�ǃ�o8ۂab+rޒ�w5�Vw�oUCD�ũ���W3����]�e�;����6���T�	A�k�T��id c1SWQǾG�k
R�܍p����=q���"�����	(�����B�L�pwn���Qn���%r4tM��E�--����d�fx��ǒƒ����fۋx��<�V����i�z`�As�H/��S�jvy�D��}�!prAtٷ�c�����8��+
~���1�wu�:�������Ԇ�h�g����oWbɹ�����J(��T H`2�u�]
�N���n�$�#_�u�G��S�D�|V$ɉ0A�.������T��<5�C�tܯ	�<7�~� Ĉ���J�׺N�b8�4��s�n��I&`�7�8�iȹY�붻�8�.7S�&<LG��zd�t㬂��gE�jA�MэP�)ℽ�UrI������'�!Q��3Ae�+eBș_�G �t;W��_r�ڕ���� ����B��*����PȒ��6z�,�k��4j/��Wd�C��+a�骑�D�X̆{���oRVi�B{9:pp�_"�X#�|5���&��w;<>���p�G=�v#�����+�~Q��	\n[��VGT�����s��>��k��Sy�s�`Z����;Mɲ�FQ4��&ڙ���!��b��/������
��T�\�Q������6~�]��E�A���0���	�T��be&\B���ԩّBx�4��g���TZߑ��*ɸ2\�_�j�cY�#x�����G��V��S��� xkU��xn⁻/y����
 :�|~��}����B *�u��}����,f'���l _<6 t�V8�bPϥ�ܘb_co���*ۄ���V]�n(��z�1r	j��������u���h���"3�O1J5ܯ.kJ�X��H��E]�6�����h���tHs�T�x���X7q/&S_�:𖌪������0D�T�q�ې��p���	țD��o��*TE;��ƥ��ߤ<w�U0"��3j53fڻ� )��)��A쬉e4��)�G��N�E�_0v�HѢ�3Ur52d���'M��Ps����%U@�	6�Q����1����P���V��8[�Ml]�.�v�*ۺ�w��3JdJ9��S��	�86"���#���O��s'��K�X���`64�J�]���ױ޿��_H�n3
I��}O-��n��A���q@��`�wݲ\	��+^��LR/�p����d��{��Pg%u���xt��`��N���4ʳk9��EZ����|�c�e��E_S@vR���V���b��~жW��F�Mi��6Z�w1�,�0>N��:G	�k�/���*�-[���Ee@D����������gvR���G��&wg�	R��!��㬜|T�����byF�R=L�֊l�U��Xj>��mNi�`�F�B�_�/�M(�{��~ �(S:�ϯ� �Te-��?(/IB�	�;H|���0��a��US����=���숴T�{��^G;���������fl� &qu�߼��,�w�����d_ ����h�aK�3OD�)�|����7NP���M����v�C���Qm�,��#��)�J�'~�i1�#����T��`X6w��ux�����)]9�?�X��%���dbm9����jd`Z��.�	�I1��M�e�gR�KTl���m�(���]��*�)4v�?��<SB	
�p\y�.9As�M�Έ�/��
�U��wu	 ��%i��Nm(����L=.�@�!-���b-̟�����ϸ�΄��	�I� �L�\��b:1��ٷ�Q�C�ʽ��m�5���NVC�,{;���j�Xf�3�'��o 
�<ؠ�LA�ȂQ �X�3v�UQD�Bw�B��.�g#�&&�\��R���̊vׅ.�����w�/ʺ��듒� p��mP(��<��;f�9�&����G�Lh���M�qF��c��6Wܽ�֤>cjH�%�I+�!��"Ͷغg�F� �2:6��,��m@���4�U)�jW۝�/�[���v�i��*�4�C�z:�fs2F��C[���DRޯ$�>V����b"S	�YR�x~����$��9���ӣ��e�W �sO߅���?�]�Ag���ٝ �e�Q����7h.Y��S�gM��Kc�ZY.�����C���)����p�H����[jY���kU/�Xwl��sM���U\���Z�fQ ��]�.�c%%�K�����M�;�+8���J{(�c��F����(�{��d�|v6W�Mq��<"�~���qB�ٖI`�vÔ�}K�Y�z�n��;Av�1��
>}	���d�-��L�����4�[��N� ���� �Wʴ�3�b3`}n	����P5�;�����Z�J������ҩ'�
ӟ�$)-OE���rR��̰, ��:һ�V�ޜ�RI�@�߽����Zh��R�a�+�:Wp!�N����jW	�I�w�xq#/�������c���ى�u��q�XU���=��\+�S��y73	FUG��l+�fe���B6�_�<c,����XKv�&\|��q�?�T�FT�!I�#���r@a��
svJ�z�s-=����˵Ga�Eo���2�9v%p���LX$�v�G�� ���=\��L�2���cpC��Wo�c�m	;�o���E�jKA��T���uȣi�1nm���p��s�K��W�=�	�l�t�!c��@���]�CC��)���m��;b�ݿ��0oOA��9