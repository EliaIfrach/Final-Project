��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
��e�����"X�iMCUa�����$w�7�B���tWEt��|�*���2��{�v�Y��Z&pG��S���̔��L�~�j.�r�|���TK|��A�R����׬su�!/��L��抒�4�}_'��9�2rƉt;�1�W�b��+܏�GڢLnd%�V�S��x)0��dr0R������߹z@oE��,X5�&�J�ume��vǕ�����|S��kwR+�\�,d�w}�a��w�5i�5~�N��Z	sD�k�]��w-=5����6��~�K<�F�o���e�~�|y0�f+*}B��e���\�>r��I�/o��2�m�
��Ë�D��<~�=V b���R2;��h���m�F���bq���j@�ӿ~��uX�_��]�8R�p��.��Nf#�bve��"Y�₢%��\j�ʍGUk���6�6-���;��?�8�棖/��NtW\ṝn�Z˳�MhG	w7bCɷ��x�-qE�\3�n���N�wIF��<2���iZ�f���o�ō�(�4�i|����2O�	�2��4�#��=b�1�m�g=��^>s�T3�|���f��yt�c(�<"	��}bt2N��鹌ԤH`�P���$�V�LO����Ĺ���w�-�Z�+�YA�M�26�J�Я���	�eh�$(� G�t��#��a8x6oj�#�d/t��ʩ�#f��ڕ�O
�ɳ�zέ6ǥP͚���2�`K�Dl��`E�{޵aKڊ�#�c�QNm�q��A�wY`�._ۚ	V��~�'b\|��X���s���-7�]���oE�;W�1iHA��(����/|-���	�E�Y��c�`˺r����BR���%�s "��\�*�)|�P(uH��gM�$��#-�E|\qj�0N�~�9-���12cAi�T��M�m2p�],"1M(�c'���Y�}CȾ[Z���v�3A4����0�,�:س60t�<?�&`'۔@�W�?��[���ɿs��i>�9��e��{>�~�^2P��9�C���sOF�--��1"��M�����ژ�-���{���εs9U�������Xثƌ�QZ�︔���<�P�\��d	��Bg?1ƱGhõ qy��klQh@����_�D�r���st|� jr?3�2�΂����o���Xt)I�Ĺ��/~M�x��L�Д�k��2��i� *�!�c�T0~��y�La�7��
4Ϋ��b��B�|U���������3A��0S:9�QYҕ\٬�.pJ�5��V]�b��V%l�u���Q�GQ9�)c�S1�d�M@gO�M��W���>Q� �-����C���f��Al�"\A)�\̹ 	DaXϡyPb��Y��Y�c�}�D��e��'��S��è���-�_����T��';��͛����v�5������^��!����g]*����wy�l�j�c����}�w��n���!r��k��G��\5Ҡ���8����qnO�V"@�2&�@��ǺL��ϰ:�o#��U�u�s�ha]ou�@�[�c��RS�_pw*1y���!RK��������0ZC-�]��0OJ��h�Qs�G�"�ȩcqs2�s�%�]ԮR�O0+�V?��
UQ�,�c�nw���{Nz�#|�EN"�^���s4���^`_R��^�.H켕W¯�mul�W�Pc4x�}#A���A��ʛw��jw�Ƒ�c	����b��s�$�+�l&��7���k��$�2�|��� �[�Q��*������f~�����R s]�E����#�c��r�'_��:9KD� x�ș{��J�T��4�K������vz 4�H��R�1Y��&�uf2c�M-�������&��"2�lT��������0�V{j��[f'�Q�w�W-��a����Ur�m�KfY?��� �r�s����.����ӂ���l�O�h�3�� 	kS�'�|x�b�ay�Tȫ�IB��n������Ot�ݍމa~8K�e�?Cy�%>�:]ܾ'�^�B�ޙ&A�|ܞ����R�-,{yo��:4�A%ΌmC�'dV�wMj�/����=�4	��4�EM!ʍ�̓ߋ޹�b�=��.�Xe7���
�^WN����(#�Gw[�Q`���Y��d<��Z9��kX��~x����[;h�@�ӷ�o>N�7�7E��pe��8(o�4�:-��M^d�W���]Hޑ��L�R�3x8��'T)�@�3[	m�H��U"�;��`)d�[g$�'�ճ�Ȅ+�j��j�YAl��
��֐���Y��Bcj�v�T\<��~����:����cZ���#�9����U@��D�p+y~p�9"9��ɤ��e��Q$.iy�޼7� ����󋬩�[���sn�ϯ��0/�	���5	ߙ�Ծ҃�SM�[�%�-�s؄�./�g����H4!l��nȣ6�8.p���Rg�x�mO��Ck���|���Z��M@�^a��?���{���<8�y�JC��}�1�a|�gh�%�OU)��D>`p�z���K������/��ۅ�%�!��v�L���5q�p��7�S�+;u)�G��˻9 p9��gF/
�`�ݍ?(�ѫ��$���ue����7�?߇Ԩ��A/b>>	9��i�a�Qp�*�F��ҧwHm��S�;�h�]1����/�{������Pm�X��O�M���a�cf�wLvcRs��e���Am��X�G��ԟ�UM:R�oy��I���ץ /�TK"��f��j#D�w��.�q����Kǈ9�dq��[h�./�Cj��X�|+1���-�D�u�,2�;�.�F���`�лvE�/�t��V&�YKS����_�e%l�+�;]>;]ʹ�!�ӑӦ�>D�ם�o3�4w����a|�n��pL9ӭ��@p%-��}��㫽5< ����l����T�A>-+��6�2F���Le�fv��)���E�D������~�`�yv<�do��1��L��=1�#�8oO�k-,�'LYȩ"��ʋ���!;�HU��6���;��]X��T}�ιϥ���8.�M�ޜ�)���<b|Ï~� �葯�|�!bU��k�7���-�s������
wdEQy�o�_��VWS%�P}D2��]�FB��1�]����q����"��U��!ᇄ��w�K���$0���X�7�f��g�Q�o�/p��Tq��/��º9��q/U5�!S��/����A�m�Ӧ��y�~A偢(8���h�_��͢�'I�ԡK.m�H��H�uF��N�'E��B�|�[n��|��}-]�+�N؍{n���Vy�x�C%��}�P�7��%�p��?���iqn��w�-a��9���	ʰ#�`I���l�W��1��S<��B�F�o�@A�v�/D^G�{�:�:�S�P�u	�����~�;"���-}˾�qw��-ً�s�H��S�ixWr`xj�ZG�A͔"�\O]�����}:�CɲU5%���J9��U�_̐k����q�w,�۴~�!����;<�����O����n��~ ��QW��<3���z*������Py]��r�X[�P�N�w�zج��w.9O�[/3��J�}&�")o��y���a���̴���<�x6�f��>������|���Xg�ݽ}:���nm&�5����mH�9)����	mw*���x�dJ1C$�
Kʧ��:�Y�&�?}�PY07��j(���Sp�y6��Hːcb cA�{�0@|w�'��Wk�8Z�ע5���)>���Yf!�x�SR�=��������[�2�I�)/�r�J��$��;<X����Wa��oaͷaw�;��<����a�����H���m��h�����֭|i�0�rc����]����.���W:�D��%�<�9��������x8y�75b>��bD�<��	#O�O��Ρ�	��6�wGV�b���B�x*RP^J���C�6�ie��:Wń�"�fB��������~LMX9擸-mGE׮E������wQE�C*�k6
� 9�\��)��t� o��ѹ��lH�?��D��Ylh��,����sՋ('����{�`<�._>�%��E�&s��hQ��׹ѥf�F��驴w��~�+�*��}�H����s�+�l�m0����"�h@�Ha���% Eǃ���'::&V�s ^}�
���b��PƆ-���\�x^�c#�3CD�#�M�B^Fg5
,�.���j�A�/
�[�k��;95m���{���S@�EK��]l����~��\�E7�I	6;�\iU���;��S�����'�J�7��~?*���: �yo��P��e����7�i�1��͊�^n�K�i�׉9vѕ�Y��������I�7k�R��S��) h�~���R�d�G��H-�Ya�n��3���u���}���BM�mb	��:��+�E<�$��|����W���;ADvTV����[� & 6��OU(��OB����;��>�>�����9;*	��#��[E�do<�Jy�H30�v��E���-c��0��#�mSק)K��F�O�W���/�rb�'P���ȉNG�|�H�vbk�Q��gE�B�8�c�y�8�)� 4pQ^�.���$�z�Q�vf[D���
���U���s��R�+pދD�*r�N��Y�b�Uu�zbā�1gb'�2���P��u���B�����!��Ԕ��O˗Ӷ��L�b"v��4�1�5�(ކd���K;-2gII�A���!D�wޫ!�����h��� ���=�3�b������������؁��Cw�1�>غk{��|-��on������kN�7�:&�|�!��^��tuN��Q1��Z"�%�Y��]�� ����}]�����L�z�sW황5Sb�v�o�l!��?�^�\�P�H�5xi������ ��vű������b̿)�~����]��<<�F��S���(��������Pَ�q�O� "�NO�6�gnUk�����@���ݝ� t�w���N/i�v݂=g]��Ȟ9���0��ʪ���V��Gz �B�����_�"�!^|�k���A.���HN�Q}��p�R��
�����a-v/c��Zh�þ-�`<�1��F���R��(N����B��@5�': �}���D�X*ЄX3��n�50�_+���b�g��pvx���'�䓕	�Ӏ.��՝�TB���2�s������5?�-7=�C��6l�Y�i_�<	���Bey�=��Ձs���D�d[Ԡ��$�doЇ � .6_��o"���r{ҽ]"׽�0�%�z�>@�a�a�+_��ƛ�f�vo�Ua�~Zx&�iD5���/B�Z�*G��p��tTx���0M�S�Ri+UkӼ ����R�U������
S�[j/��*O�AV2L���ƨe��S�3�ܨ'��ł��0�,�o;�^+�]M�k?�2V���LfAmm��lֺ���GA=�^��*GHO��A� ̖�:�>5�m��̚�y�|k�q��\�6�J�A\q̿��6ר��Y"٨�N�+��[p0S\u¤ﻈT=Ӡ�s�&r�
4�k�3���O_1���gmB�^Ʃ=��%[�!N�h.CQ^�FQV�K)�;��t~�kЁ]��ImN4�w�/�k�u��PѴ�>���x�]9���|��"8onM�tw�9��C;
z����\���ɫPXʋ�D@��L:�T�L5��i>0���i<���
 ����̟�
CMh��)�X�:<�J�ٓג�]��װEךD�B�D=���ѻ�!~�X��l�m�DR����RI$�O��Ӕ�d�=&�0�����|)$G���������~yN�<Y��u�2L�.��Q��L��قI�ﱐC@\���$�u�}�}|c�I-����
d�Qx�؀�ف)���3 ����n�(�3%O��c�'��?<�^~��n ���Y�xv*�κ"m�7>���O�	��X	�P��:���C���/Eq�<~V�L04�%�ZY��s�,�t?5M�^*�s�Z^V14`����8[�ob�֛�i�svޣ��.FKj�h⢜�xּb8kή��Ě;���̪3��e����`�%�/F��7LC�qd0���	̙��4���Q�5�a~���{3wՋ� �^���}�K�{�w�6�����ө�� U�:X�Yc�)��x�A��9���#|���3��G����ᓟ�ݿ�p_��z��OR�"�gv��^��`.�s
��\�$t�)������5�=0�������r?���ږ�Oq&�]��CpPX��[��-iU��Ѻ��.
��KA
����QF����q ��'�'�/,#B���?
�~3�-d��ߣ�������=J^�Aw�{a��u<]�O�F�Y`@��,�@�Ϥf�q�z���	� k ��7��#�b|5F䱵,.S��[cw'�N���{���gӞ��B���Fƶo����+X��(ms�`СXc�?q��;�eG��v�`�E���L�1	�l�n��7R8���?uX�V'we��Ҭ]*��G*�a����kb���@R�z�Q�P����{謫�����=��2�p�xWH�%ZT���ދTB��h��$1���G�i������߀ʦELe���O�[{T#IVuFv����'�@�.���AaVN�.&�6�[���Η���3쩁�Β�.�jJZלyw�z>��"�:�1��3qg�I��rBj�r}��(J��6Z/���t�-]�7��g��% ;69\�i�cl�l�`� DM��Dv�g�����e��f�H���EJ�iy<��K	�.5QGҵU��B�wMr��_S�Ӻ��f|>2_�|((�#�4|�!xh�6|����s1n"TB)���S����Sߊ�z�e`K?V#��"����}����r=P�@W�eJx�6
���w��R����2X�}Ռu���Ac���%|�*�tG�3j�`;Ǜj�}�*�����zح�X4½Y������㲍���Ԇ��W�(�U�	��C�[ʣ��2�5���i����A���r� �H��|SDϾ�ۊo�x��"Q���Ǿ��*�M"�C�^SH����e�w/��z �㬁犐�`n
��?��p�QU����� �K͍D�-,h��8GW�����5�-dߊ#���K���[��G��з�L[��~�0���B�����tޛEӣYZ�^�-h|�k�M�3L�1Wv��ШGeV�ȃ{�"��U��S���ڄ�_8��Pd��,���{����Q�~�SN�[#y�B�y;!ƚ~2��J+!���������Nf� +Ȇ��7х������r����>�~���[d�!�@�;U���bc�Z�&�>�?�}�?ZʍG�EQ}ѹ�(:!�>`��.{ހ����w�z�s��S%*� �O(<&�t6�7uT{����Ŀ޳�����Ȭ�~�Q>}�O7K�X���$�\���L�e�����&�=	J�����Wa$ FrҬ�<��}�8�P���
�̮P�~����sd2�NzKǍ�Z1�i�w;��(M�NZ��,��Ү�WzO��eɡ�ix4�^U����ˈ	�=j�-��G���IZ�F�EX��dy?�S�/��1:�	Aԉ�BWWb�1��ͻ�+���γ�$�r�o�QOx ���O_�ʄYo���aW WzfD��7y�:�畝TB�Ff�k�����]����M=��T׀C|/��R����#�j[{�MH�|��>�ҽ��8V7�F��E�����*�-��4�!\��v<��E;�^�+D�{�2ax''w�?��Ƴ�h�����(��Fc��T,Qkx>?:H�}"V�l��Z�8l�yԞ�H����ʴ &�<��$�S�/?��r��o�DX��4�%�&��\�E������Я����֕�|䳾1��khe��9���O'ep��4n�i���e9�>f�qN��'4oM���f@�p-������Ŵ�(17FC�BW�lA�#`����ŬUdVuI��7�G�Ǌ�0�	�)�{z�^��\{j;8v)���@P����ؒL%�"?Q�G�2˱�!��3q��S��ޛ��G�Z@�7x������أ�r'��;��6cHmrٴKح�Rf 0�����z9�f���;:��dFo���W�K#�qɂILĘl���=$�cRl,H'6\%�lH������]`��Hl����S2P!V"��eXEf���\\[0:7ܫ�3Ց_�|�DH��b4�)�^ h����t��p�S�j��4Ѣ��o|�!�݂��h�XKb���}���BaW�y
��)[��JD3솬������e8܃�n�B}�e��J��pЅXI~�"�uSl�ћ>gl�nƑ"��c����A�]#�ur�8�x���H�(�v٬��?3��!���	̤9����t6#L^a��ql}d��Q-/`z�13(�根c=���j�z�.���b�U��˓1��,
���>U��a�=�s��2J���	���V��?M��X~Zd���%'6�V!����b�zD~q�Ȉ�d׬���q��[h*AҒ��ݴ��5�'���ey���-��<y�{��\g��L�)�b�C�镽�{��g��(^:Λ�EDy��+���r�?�-N�$В���rn˜��� �^2Z^)�ꃇA!�G��UH��e�t<�	�VyÔp�i�6� ��VK�͂���Z��Vt�TM@���ޱ˄��du֭�?��O"�U{������<��JR�O�1�{�S�"�"������J��������N�Cᄡ���l��P:�.�˓�̚��:��X� ����p=#ݭ���<��Wռ1������~�0[�ƆS'��1�D@L�Bq��)C�Ac��)gW�2���@���
U�#A�B7&�f,~������xg�B�ꏎL����"�)�v�� x<�{zk���z�A������#:�u�lۣ�ٝN���7�^�:��q�B�@�6dr�`m���Eo�ۃr<^�HRp�[�� x���P2�W�c�2����l�5�S�ԁ�����1�	� �qEA'�#��ظհ�e��Mih�`$ �=&M��F)�oM�s^$��i�<�H���K!�ϊĥ!4%��٬�Ao�{�A���SГ�h���F� S
�f�G��w�/McR��\�~�~��Q�ꎇp���w��r�]t�{sn���`�Z��~�j���c�L	��-��V��}K%l�8���>B�Z�� v٤�l���/6����4�Ģ���f��<Ex�O�쇹������c�aX�m�z*�1v��5�R^�k�������Ӹ�:!�� ���� �Å�������L��:ņ<�ӵԩX�J��,����Lu��$7g���#;�*�FF�-�*�I
!"�c��������;?��O����]����BԢ 
�=#������W��`�/
[��y�%0���m���wk%8'ˬpw]�]�	��?��"w'�&�r��ӽ;x����2����y���I��)�j0��6��S��g9��*�3[J��y�@�(���Ed^1ME��(��������r���@)�^Q�1nLc��X���XՈ���6찃�#�ߗ+-��������C�U21M� 
��E��S�:���B�(� 4����S�']�3�.i�HR��Soz����ʰ ϶_��/5�D-�����T�Xݱ.�\y̺��G�j�N��������f�����;c(Ѥ��y�t��
�,�BH1y��|����D������t��;�Qbj��}�}�A�h�V�$���ҫxFٛ�'�D���o6�x�Gy��o` �+�1�(�_�5%'Ex�g�V���'�-_O���t�ǣ|�	B2����A�Х[6g�My���k=�?�S|>
��ǈ���*/�n�,�9�>Y-�혗�$*qєŕ15�.PRy�줴'�Q4w�	A/��,��T��ȃ^��{%�XH^�)�Z^�1g�N3.M�n�]Uo���tէ	oN�,
N����m����#�x��oZ`o�B��Hx��:DS��] ��g�<���ʼUk�m�I�=�Ԩp}�Y�4��AG�J���H��d��y/������An�z�)6�|h+�@W7값�`x^z팒��^o j	W�푍j)�,�y,|*P��KY��'V� ���/�tlV��F��0S
�[��V����!3�R�(�(!xKx%Ȗ-�I����7�B�I����E�"F�W������ܕ9n~���}p��� q@w�I�5��2��������/�Ș4 \*�X�m�<,���^��/bh.��ۊJ��l$���*��a�ouHz�stT_I�����5�%��+^����P�i|�3�s�ɉ���+�!�1����H�}�5^�g��b�~l�:ڑ��������v�?��`��� S6Ϲ�@A���������g����a�H�eY���i�����z�ٟЋ7���m_�!�f^�጗Yz�iL�8�k5d���[�
���6Nc�޿�*��ɝ�4�kI|��O5�
���w���\m��bˏ�F�>,W����@%�e���7�W[�"��e#� ��kh
2����(����"���!6̤`�o8���K�������TZ�@ॹx뽰�1����|o7@I����hn�./�(�M������c��Lgu��5�)��N".���}fQ�
C���Ο�i.V&'�ƻȯq�s5�[Pb�1�D�T�WK~���Y�#����� �sC�
ʷH�h�:�f�/����b�!Dv��Ԏ˟��m��#L����Ҧ Of�a�&���� ��X�􀎽Z���j c���Of�a�@��*5+/���n3����x=,�nu�;	1��XGßN�ix,�SB�����E�y¤�r�A����~%�9���3��pR$���^,�?�J�l��ƴsxxGo�o��\�R��s�¹ظG�h<�A�Mչ�et�8��3�𝁽˭���g�$ �K�BӟUô'b~���2�~�X�� J^̪f}1�~�2K�'�O� ZznF�$I�sa�0�.�!c��8S�(%���!2
�r��W�z��wR�c��m�/Z��=���m3=�RY��7�����!b*�Z����W&�L5�s��-ϤX0�!����>'����9�
#��=}:/����Q=�K/�v���89���6�ӟ3�@�!mDd���i
��}�QQg�3�!�r��)�>�2��v����`��C8�_��,1� �t�_/�x�������2���a$M�W$r�����4ZN�m���<ޭ��W��I7��fQ�
���#��KAܙv?��-7[�;����'��V�S��.E!A�+�v�YsAQ��),�I��l�I(N��H蹅urV���4��>�L�J�>�Q�t��<1~�,I|L>�æ�s�>�>����*z62��:`���Vp��7/tPcJ�3��Ղ��F�ɑ�t�O'r��@pLI�Z��8�7@.nI��7�F�1w9�J}v���a*�[�w���0eP��t�����>ơgq<4����l�R�@�$�ϩ ��Y�{�gM���ў�*6@��^g|�����K��2r�?@Ѷ��U/�� �o�H>��xn����7i�Fː1��S���J7[�G�@nkz̼N���`�y�B����<pw6�L�mz�[��=��i�F&��^�L$�����"�sP����:��s��p��yï+%��]�&�Fئȶ�,��(!Xf������R	�o	,:���Vp�Q%��J�4�,��\��[İp�NB1y�h>?�h�ђ��MX��r���)?�iE϶rW�h\Yfv[��w�N�%��\�*kBxA���D�@��,i�́.��c��WVӞ^���Z�wFJ8���\�m�C��㱞ǲd�o+���J��,}��Ža���
'���>�t���Y��$��٫��m�L�(���&�ڡ`��1!��* n�mvHR�N0�"(����j4HF^�&P+��9cr��Qf�`�F+��$��#j?]��Aj0�:�*[�Y��7r�*��:��xȝľ|HS�y��R����dfԋ=��X0�0N�B)c`B���O��~�кДR���YX���t�s�Xe/�'*cn�3Z��I�o	��m�m�	����6�2�H�T�A����m��~*�>�u���g�4S�Yqtͷ��^g�2�����bO����!��Zz.����(�:Z-⋘�Ze����~��O�|:pF9��Ԏo�>�S�ݛn�1c�pd4-��"sd¨��؅��B��@;pLs]��SVq��Bf7O�(�ʚA����;�h��c�q���T���e����y�0�`M��Ϗ���$�몎�y:瀬��?��T�k��M�3z��� Ⱦ3�ȳ�&���, 
�%����$#�ΪmO#^��"NjYAԈEЙ���2�����U#xstbkv�������n��m�z=zg~S��F�p�<�-C��C��;^����K�fVY����&���l�q���ݶ�m_@��@؋}D�/��#��̩��f^꾼v)�sH�d�p<��b�3sX��!�u��?H܉��$̊Z=��[�<��4
!��QK�Չp��EDz��kA�5�Ĳ�ӡ-?
Fʩp�w��4�W��s;(�c��OXFMh:Rz����NCt{�	@�V��&i�mNu2��2L��+��f(Ͳ��(����B�`7��b���Q+��ͤ@ȟ:J��9���Ι��z.��RjD����xpL��̾��I���e�u��Ɍ��9w3T�Y���}����f{QL�b�֭��A�9����T˹��K�J��cyΑ��#<_�@�Aqs�X�*�����+�� )���V
���U\7�ʋ�j���ݺ5�ɕ���#4�Ɍ�ё"��_G[�>$\���_�i�z�e� ;B7�G���W˕�f$MT�P�nW�aM]q"�I�$�0w�"�d��lM���i9�W�)}K��]%w^FU�����`͒��~�e�!�Dޖ�UW������/����`��B�����
Hu��9��h��BY�}3h�-��I�u��C��K2|��:&�m����gt� I��M�[Y7U�61[N�G�O��:e�k��F, %�C�պ��-�1Χ�1o� �B|=�y1��E�>�<��T���8��l�(`16�T�|��5�ZgF��G�?'C�^�j���Cm���ys�C�Ĳ�a�K¹��0���W�/u[B��m�i1o���Sk蓙����5�{�S~�M�q_�֓�5��	�$Q}o)bk�s��?�����
� �����Ik��4�bY[R�&y�C��X�c���Czh=���'a�� �������F��$	��a)���FRq:*A��@�ϯ�,2����յ�������j�6��!��Bz���&~H�m�l½�'sY'��[h�<�G�&S/`���fte�r�սW��^���u�m���;� ����}Miq|�f���c��2�FG�56�K!Z_��)#B�`zz؜0�ˠ|�1x�:�(���M�E�Y D�Q/�M�M�R�����Onja�}�5U�C���N��
��Y'�n ��E6*�� ���t�:B���Z��=��D@��l����rH$D��"�G8I��.�Y٫���Mݥ�oh�������mS������."�ŉO�Zr��&�ƌ�dj ���XuڵMc��>Liֲ�S�n�ˮh�"{�#bij�����N��6fٜ�N篶�d*k��K;٩9>IV��� ��z��=��(�] ����v�x��mN�L� CyZ�l~�������wL�,�0��Z����=��;��� �ܼ�C ��8Lc�s>U���*R��9I/Օqt)O�wb��߁Ԏ������=�[�-;j�"�D�%�Cb�S:w)`'�1Kʲ��_]@��C=t�6�ư��1�xNT�c�I7ԄK�Њ�ɗ&�K�"͋sw�hB_�Mޚᑝ���j�=�ױ�9^�I�5�D�ߡL}|���&f�lTQ�zˬ&ۻ�*{z1l������Za�~��U}9+���	@�CY�0���8L������D}�CpC�(^(BN�,.��Sii�������w8�fp��[��P>���ǟlxm��0\��(f�~҈6{:�L�J+i��(F6^��V��U��.1�8âϵ���T\��<���@��0O�'9�@���#5VӍ�n��]цs+��~��QfE��k?�ۋ�U��*C�;sm�2p�h������o�Aۑ%#��ui��g'��(�F�K]�xv�3��p9V���G�,֎{Y?��՗7|��n%�֝�blA�C5�4�����)o_TZ�j$FD��T��x<M�X#~b�s��Z��VSocs}P� �!4��,?�4�l~�\�R�V'�mw��Ϙq�z��r�b�͐�f!p(���+����<
��	�[�?pZq�h.�?g�^�z=H�/�[�.k}��O`����D=�ħ3
����Ĝ��ۃb��œ��� �a3�:D���ZtL���z �j�
�w�E�m��4j���o�1'��6;tR��%@��������p�&#1��BWk��(���7�1��m�����%��Un���)u*�T��! �Io���*y��]��gQ>��91��C����;��!��']~|E�ьr\T��5���#���pY,������)3M騛Ѽ�D�jw�	$�
*�HێU ��&1�4!��,�����B$��@^�D�����j۹��� �Mg��Z�����dZ�9fpA����Ř�Ɛ���#��J�����no.)8d���􎻣HNX��E���[���O��ӽaM\頍����9>.q�i~���9�=�tB�냇Kun����_�t����	������ⓆB�ԍ��s�K�Q+W�ّ��Ą�n�i�N�9�i�(��O����̱j&��ǀ���"��~,��������>@J��Rߓ,���Ѭ庮�T,Syܹ�)>�[S���<���x�
�M������{)�졮	ú�)�R�J�����E8�S2����;?6�u�_yd5Y/u�A�
3��ͽׇ/� D��s�ۑX�Gչ�3't���G�bb���.?a_@��bG6Wj�tB�"��z�E.��͓xe�j{\+XY>��|>
�:��N6��&֑?!	������G��N>� ���'>?m�'��x����$M���,�F�<~^n"	�����I'9�+>�Y9ܭ��9�I�8��ݴ�i7�j�sz�c��%�������^�ߥr�0P@�����[�V��B���D��?��5	����w;���셢�5���ssD��K(!�ᘟ�d-�d�gx�[-�b�*ZƖ��M��˩++��ݼVjG�$C��/A|q�<�t��uN��l��k�Q�/�|'nY����p�&J:yl����2I�0�qP�J	R���ԣ���&�FI�c�d�z���?�%�	�	Ʌ���d7�XI�SΠFSz��)���L+o|[w��{UI�.�&/YE���]A�W����V��!�'ʨ�2��L
��R����k}h��֊�zd�N�T���P�=�!	��?~M�΢�`04�е!%��
��>4A#1��F݉���(v����Ǔ5 8��iǧ��!�aP�3�M�^�\��Z^<V(��J�}�����$��T3j�~�p����2X������/>�`n%��|�b�� ��uW�d�Y�{d,8�`�=N�G�L�M��;f=in8N,`vb�Zaȉ��������3��`$$��
�h��|�����yX���ຑW��p�Йj3��b�d]ou�
S����+\���T�����b�Y�l�z�(A�ߘ>���]ҴX|�߂��ue��^a���Nxe7��"�sJ���8����w#0S�6+�e��m|��>A� .`}�y�y���� �.m��y��I�~G�z8����$���0u�|pƷԢ�6��;N�Ȯ��i����Xȋ �r]19�	,��-m�=���k���_��	
O���V��?՚0� V�^��b�BQ�~~m)�kR[҄b+~ӥmܕӨ"��O����C��U>An	�m��S��$:ONBؖ��-��& �cdT�y��o�JJ
.���_l�gSC�ߒ����(i���6F	�%������
�ڡ��rh2��9��H*����*w3��ϣ��W<ji�ܬ�%��r�UGHP7/�-���{�ge�e�]�W�����r%�|�,���5=��{`r�����3���N��&;������Mdϋ �C�v5����>T�ǲ�� �ġ�M9c��i���m�9up����fs*!qN�l�F��C`.Afh Ԟ���^�J�C{��ţ�z�8�h����_����ɋ��Ld�}����
s�y�

�[k�����G�|�e�黷N����� ȍ���KY��6�O��)k��g�Vy�_h����%��'<BYAg"C�<q�=�! t��CK!_�\,1.���8�v2�C�˕&}�E� C�.I��(�q3�P�0�`Jm�uZ�Ř���'�@�ĝ�K*�ǁ��y����5�m��&��!�#��W���R�!�$�D�"�-�-2l!定�4d�s��4�qn:�{��HL
��O�Y���]�ސob'��Fc�E� ��v�g�(��?������W�_�%pm�I����X6�NM���ڑ5F0D(�@��RQR����n3�U��3�W��?T�"Ϗ��o;�w�X��G\�Q%��aN����j�T�$O�3zv���=�Q���?��sF�<���]ż&j$�k}�����@@S�&�f �%"��:��\��_<�5FL
�5��[м�4*$�lg�%���"��tz�L�dO�َ(�Y�J1����g3��V��R��{�b̼`�jڽ���S�J�Z	D#����|O���>D��zt����Z�8�F����L+S�_�#o:R�6�~��Q����񗟿N�'�;���.y�ONҬ�z5�H�6�)�Ӹ����u3[���'�U��p�ZX7%�{���z_^O`Ay(���QO2߳�^��U��`�(U����E�?��3p�O�sV��Ӝ!�m)���ZPLm�{6�7���4�k̀Ac����3� }��@ʚ���K��pM��T�6��)���W]1�|���1���7�*"�`X��R�:w~cYt�2��<7�������WbT�&E�/۩wt14�4�è���p������	�6��^���oǏ�XHBԬ��ˇ ��)�E�̌`����
k���# ޱF�f �_�����|��K�a;��oJ���(Ě�>��g��"�p���+��̄�K�y�M����:t�)�O�F2�Ю�������Fa������5�k D'�v���k�~�/3����%��oph#0�ŭ�r-��C����{X���yvS#�����)
����!B}w&�fe��a�Ǎ1�/ow[{i�>P�O���t��h���|Gr{i!^]���z���ٜ�}�j��M
x��'���G9�Cya�t����|Ξi�{�]߯����ɏ2��,���S��;K<����RUA����D��fum_�l6b\A&}����y��f�����lh�}m8J�s7>�����N������~�4��v!Fј�AXN��"S�N4BǦ_@�� 6�?:]Jr4���wߊ��9��k��Y��Ľ}�T��H��+ݚ�F?Չ]zy�OGYb���U�A�ʍ��݌�E��z��4Rl.��VkPeH��ֳN��ƈ��'��3b`���m� _"$#����P*�P��^�0�"���i��Vr5���S�d�}|l�#����q�}�->n�ı�t�|�Ԗ��M�#?\f��?,i��"��R����m�˃3��ˣ�E,Oz6X� ���,�uP��-&��/�
 �P�E`�ό�s[86�[K�K򴿬�9�
��nqb�� Z���ӣ������!���ȃ�2w��B�K� ���:`�H:�KF*��݇_�z�r��Ж��6d�͔����H8���b�'5��&YF�/w����/��G�c�	����a\H�[|�}8Yu!@y���B뜒�m�␒��"�L��7"��T"�i��Hv�*?r1o��a�S�d�dq[�
<��l��I�>�#v�=gN'������@�ګ���V�qV���nR���s&���5���M.��+�	^h�y7S nU�O�6��:(���ߟ��y��������jf�4���Q�z��e�d�<�-0�+�+��*�=�C&e�/y�-��O�pK���5��X��W��h�R��/�."(��O\�xQy������9A)��R�(FA�;+� kL5�gE9���D�Q��u֊8a�h�D��X�3�������χ,e~�bcj����X��@�A��!P�����z���Ou�ɝH{3�Vٵ��-Y�Q�DQ�ЇK�M�Yʳ�h�s�����n�#�߳S��7ؗ��\�_����{|�x������A��n=�:��Ù�rQ��(�5L1oD9X&�i~�^'�'��. �aaL������`(On��gVv�<'G�3@������R�~��/x\��K-4�($tt�I����iQ��A�]���a�bDb��d����K�o���7(���~���˟��t�X_�;�!�^�6,ݷ�<ճ��H�m����wPƁ�sU	u��"1f���e��v�'xψ�Ky�R�Oi��#xG�s�����޶�XD�Ǆl9�`�yή��V�%���y$p-���Fi�g��y��ͥ4Y���ؕ�6@��vZ��]����>bݯ��(�miۮ,��d���BG�Hk*�\��П@�z�@�vJ�f�T���p��ԃ�� Y�+hOv�5Xɉo��7d~�q[��γo	��yq �`3Z}���:��TdI�z<N��l&�a~?��WU�f���{qM�/���}����6X���%��Z�!92FVA�;6]��{�G�=�##�sB�'�d&	�x��)����	om6s��xKN���ܞ��=2��n � a�p�ՙ:Q��Mt^�)l��5�.���1�M��͓�?u��g�h�S�܃�aVG���W������p^1fҭ �z�P�'ac.���]���1�H����4���h�V�w�Q��H�����[X�A�oQ���j��x	�:fS�%�J��1[�
���2��Ht�<6 ����'����/�x��"�7у��J3Z���/OB��*�c6���%r�ِ�eA.�,�2��y(q�}j�&�P�5��u�F�y:��2�!7^�@�r�d�q�Ю�����[e;���5�HZJD '��Z�0n��_\f��:� uO�pN��P���oF$��N{�E�3@���&����I`pl�
F����b���̏o
�ܳP����>)����ϵ��]�b�)}��d�
%�J�"�\��
E��<�#Ϫ_�%���/��z�P�R65�m����uسfc ��0^7��(�F�����=g%��}���S���[ũ$Θ�6�U�ձ�&�H�xޜ����z7�L�Jm�{�Qpau��g<X��n��>�΅��HS�٦����T��f�����H�b˫\�t:�����dx.�H<�$�7=jD�S*F>i�
�J�w��Nz�[l�ϳ$�<�a��j�(�6���踔B$���?U9֥�[Z��/�"�*��=��"��D�_$��ր�Z<����0�����<�3xI��ZL�)�荘f%g�d&yɝ%�T�Eȹ�����L?ж����Y#Gwg	�B�����HX�{̦RWG���rQS�V?r!�s�;�����q��H6�T�hg����7_�	�@�3Ɯa��&	n_jz@�&c.2n&R����zQ�\u�C�`����"�͒����zJNq�)!Ǖsz�>(�ʴ�]j�Wp�+̔����LH�9cn��͓a���rgn�!�EM���j��!x�&t8`�t�zp���#���b�t�gS��
�A	d�i͑�{�����t\�+�Ct6����!���G�D'g���������|ϒ Ѐa�?l@Ȃ0�� [���_s.��p�h	ϕ�Y�T-�F�cB�K'�'�p6�3V�m�t����KU�,��Fc�j����#-ޛRi��?�sS1sE����%�U�1�$�Ln�vu�~Y��8���|�Ll��fJOe].]C��#�GP�t�M�X�x.Rٽ�!��{i�����ܴ��_��aw��7�(z	S���B���|MZ��'
�fNhoc�j;�ͺ�y�3Ǐŋ^(4?�k�pr]��s�h���]����(9߁:X:��:MN��]%��F��R�"�5��-]���j�BE���>y3�����_#^�ҠwE�B�m��<&g#�.�;:�k�7�џ�늘�ѐi�b���)/ɿ�$W��_c�>��}$ok��=>dWT��mM���i�[��&���(� 1�*#�UB��O3��+��#�E9��y��ڲB���~�VE�2R}��F"�8�eE7J�=���r��h��<�2�pm��r�b~5���]�vdx:������D�Q�yL�X��`�۟�,�.Zr1ԡ�A�#��� ܒ:e��Q�ݶ�^r=���&��R#fg6�	H v�Y�|�f��~��=�u�Zi��*�N�S<?���/�Ӧ�ҋ�
�Zal�3������Б2�M��>���;l��!�v���r��)�Ԟ��(m���J`m_��ٖ�i؈�\�藴:�|�t�h=Rt6y�6K��B���/�7ʣd��$D�5C	�fb���R�kY����?����6�ng.q�:�%��}z�+ɔ��"rUE� �!T�ؤ��Lܜ��A��D�s�4�D���!�n���Y�����|JX�t�ǳ�"V�>����SI��j8X�d��dꡙ!+�\��|Dy���u�xn$U�<��I�$.�z (�0�E���i
�TQ�ҿ��`��zt2��;=i�4�R�t�/�!���0]����X�!}�cn)���T9��yx4Dx+[��*'&E���X����(QB��i6=�$�k���Ж�=�J�TuQ����W�w5?���9�益����q^�5^�7�Zy���
lkP6�ʌWW�����6ךpa�v�sC���?��nCMc]�j��q�S�*��5������2't7���|\�x�6��n����W����Gv�+�5�H^&�V�Š�j�Ve\Ao{VaE���1��D�Tft��@��L�H*6@��cg��ﴺ����Q>U��x"T��C�I-x�& �#0��ӕ)A)RƧ(��'�\8�e��
/�Ft�-��j��Ay���T��!Yr�fi�z	_\����cX!1a3*YN��:g�_�l�|,�hΖ��� ��K}�w�z�7�_��vJ����1��BNv�U�r�#}�{�k���s��l�9�]�	V�{���w:H�Bt��l����:i>��i�Ǝ<��VgG���O��^����\��ձ{�de��=�N����:�I�r�7v*q�7�[���k����v%F��	��':`��t(��@��F=d\h�	�����L��<�,����ߚK.�Z.�A��8`|ϸ��h��"<�Tx�H��ķkR�q�p�{q0O�;����D^�@���Z@'�wx��G���\Л��ю�M�;����w_��Vܦ��h����[������}�(خ�R�N�(�����,L�L:�c(������u*��+��d�H�SI�E�Zzm�R�z��/���3�S>��bZ���	׌4q,���j�$���Z�@�QW�mfY+	�N�����R+��a���P�͏B��me���,x�3��Ej��I�ciU�`=�$�8K%<i���迗3�Y���+�L[K�Gu�F��9�vl�PqW� u���=�DyN6l�˧>�ɤ9�b�~N�QD�41�p�gT���}	L��y�MFc{�\+RF�DR��8'L�|y�`T۱
D���P����P��_h[��W�v��d=N&����C�c<u�̠�s��.�E"���3��83��y?��H����ֿ%�QP�@f��2�3�oEWWI�Y֪���ʶ~-����������͎T?
{o�������7Q�#}�ݥ+N�#��d�u�Y�x�<pߖ�j���4lqb�������Wҁ��Re�7Aǡ�C,']�n���q���N4s�"��} �#�(2�ˆ �B�~e�UD��V�`���t9�E���a��Ù��n�x�1�翽�x��P=���.���_�f,�o��]!�Kr��c���������!��&�Xh��9p5���A�[�I�N2�ZIC��j����#��L;��L�[�p����(�Ԣ�bD/�nh�v���u��YP.0{���`,�"F<���a	�{�+�a�|m=�eY�y�@�q4޼�����^;8��γ@g�,��������l/"�%�p���f�e
��k��ʳ�ٱ�5l���@g�ͳu~�Ev����J\;�=��E���'K��c\K��(�\P@ef _����)�iVE>�YA�Quq��2���AmS�l��t��
΋�f��% L���*:Xq�)�X�l��^ �;,��"�$d�`	�9��#s�6r����$%V2�ܫ��k�Q�XDa�>h������`���m�Ɇ�t,Z���~�59���i�~�e_�	W��5�g�3�����7&JNB:���8�����3��#P|4��g[wT`��NvBMkQn�@J�6��V`�m)���[�k�y.��-�P}���%��~_~4��"]�~Ly�Kj�)0J��J��C�g�g/��=4M�"B��W��HJ,0��ط�`ϵ`�a�[����j��тD��Ή̧�GN�g�5J�t�L�f�����i�~ܟ'���;�LL��f����Q��~i<�,����Ԃ�4-���zOu��:�`^S5�oWhM���^��#���f����xC�ŀ�