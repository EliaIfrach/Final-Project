��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��33�z_�`�f����EW^7"q5���K��Ҋ���CU���w����=G&�ʉ״Tĕh�{%�E��ڀn[ɥ�'S0abx/���s��n�	�R}��E���n��Oq�9��>�\@����?�g~�*�s���}���X��#�~���U"�,�'�v�}ks&�iK�K�"�����0}�6꺍�}]^5�c����g�A�v��}���d{}|������7HW�!wV �Sn�fdo,9`F9�%QlH:CQ�p�!DM�5�6�my+�<M�~|�\�o�@��b��E�Ë�$���央�?�d�><����=·գ^���-�L{_3:��ُaK7���$���)zD)bo���<�m!>h�nW��6���ɯ�d��`�9ƀ�#qK�캅|�����v��s��C�"���6�0:z��D�5�m�̻bk_3J�U�lm05!��4WR
�i��"�=�{<� (~�Ӥ��E��U��� ����ٱ��j����|�c��)<p���rԯ��d�0��Ӑ�:�tr�!�D�D�M�G6���㍢��v <���Z����1U-��۩��F�k�Cdɇ�@�-�ޟ�e>�he1�(���vV�΂M��Cv�}{641�7�6���u�E����o�*§	-,0�u)ɍ�'�6����7�����A~��(S/�ͱ8\i��/�}�7@>y��Z�h��������:?�CɌ�#^��Ɯ��oƣyr��=���T�	��08�W1���LWc�a̔M>��t�-�)�Z�sA2T4=����+���Q��X~��U��!��+ț]��H_����jR;!������ԣb.�{/�x�ΰs�k�%�f�8h�����aGT�D���N����ؑ�T\jSFփ���������p����2f�	��_K�C�6�2��<���[��|�٥"ݣo���.�"��E҂�e����`F��&�wU�T�F�]�`�lsDm�%����X������������Q��*@�_0�y��uױ'�A��oM�y/���?q�[��Nݞ���]�gzS�!���JMh��/>��M�zU��J�ܴ$��v���×����'t�m��Z&�9,�
��� l@���@+�;�p]=�&9���g+c��Θ�U�F�G������H6�Z�U`s���6+-ȲM��������<�I/!q�U��ˣ��{�9O�?�ډ�T�2�%�*���{����S�����xD���kx4R]�lU�2�n%к��M�M^���=�'?��U{(L�jK}II�)�lVZ����e/�n�;O�%��dsK?>�#�~R����
�ct�n�z����~4��f `Y���Lə��>q3���I��}�7�<�I�����3-hsҠyM�潗��i#������;��ISj\�}k�=v��%��ʗ�gɆ�7m��y��+T�yU�xg��)�3u�md����T	�4�'��<��yė�>ឥ��5x0���z[۶4�:\qm�$Dc%�&��N�\��9"C�"]q潶����ƙ@��)K�0������}��Mg�L��5≣�� ���C%	`ʋ���^���׷h����Lg�����w��&���{3k�<vjp����i��H���<3����i�D�W��U�N��f�S$8:ò|FPɐx4怋�5=���ݖM#�
4jv�{�����Ӱ�y`K���L軛���ǌ�E,��P� ײ��5�*U�;�R�_�ӛ��n=TF�T����iD��ԝ{w=�����,��
�+4
gr��c�{2I�Ƨ��֌¬}3J�C셠~A���-<ʧ��%t9��'k�Ы#V�#Tl�&�����2��C��|�ro�n��µ'_��m
`���=7Rb���/po�.��nf�D�_���oC;�qpď4�\�����R�HDD&��Q�.�W�s�o��
��iUj&`99��|8�����CP�GL�`Q�+w8��#�`(c��-�G�y���d߳��mN�8��Su�[�4����W%F�����?T����xT���`�.��H����6�����Q+�j�z��5�W��"ᢧ|ɸ=�ml�cb�S�	����L��^��1-�� �%�����b8,��# O������D.#w��U}7?=/�ɂ5GTM��aZz��W�a�cQ$
�yg��<���<I��;Da��,S���IiCG��>�׺*��i�%��G�����c$ğ��$m�L�Ϸm(D5A>���y���j�*mWFVT�x�mc)U�����X	)~���IS�H�ҴUa�T&+�Xnc^�{<eW�N�N��\)��~�,�n��a�c!N_�%T�:&�ՄT�]B�ɦ�(��w���%;�D6	�x�D5,�W�qB�0�)i��rvE\ L����o�-��?u���J��_�Qgz\ZI2�6	 tR��F�%?B�㌅������������,� 6-��̱���_��Ơ=��&���#�$p�s�����Hy;�ψƏ����Ը��Y+��!/G��I���n� ��%��F�S),�o���b*
��c���q�^dWY��<?+�Z/���@�]*�4�)>tkI:mI� f�4%�j��3�n!L��X6�0}�"��q9 |�̝R(�{õ�3�D��Z�i��E\������A=C���c4�q�ٳ$6��p�ڒ}�l����BZ�j�`՞>�Ca�;������m�d�'��v� @�2�M���6Q^�w�������ez�����$��L�6���X$�x��A�<qG l��Γ!�"a �BVK���.@]��n�q�"#��&,Z�U|i�'�� {����M|ʺ�堉2?4F=�Lk|� ��w�ڴY����G� h����	�g���d��PHm,����K�"����q�R�d�@%*��	ڎ���Ha����n���
��5%�A��OKr*�z.�eXO\��H ���sF�E���#���)�"�M`SΎ���\[� Pt��Hia%ĝ����3-����c��K�] I�d���� Uz��g��uǪ�6�� �~bf�EΧq��������1�k����!I��Wxu��[:�t7�� o��9�l۰h�b66�ʪ�3��-���PQ��}��Nr4���lК������*Z>����bv�i��9Xt�]hJ�G;T�_���`q��mIy��a