��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��33�z_�`�f����EW^7"q5���K��Ҋ���CU���w����=G&�ʉ״Tĕh�{%�E��ڀn[ɥ�'S0abx/���s��n�	�R}��E���n��Oq�9��>�\@����?�g~�*�s���}���X��#�~���U"�,�'�v�}ks&�iK�K�"�����0}�6꺍�}]^5�c���@��p��� ʂ�P�w8yTᮏn���;�l[?[����a*v`���ƺ�^o����l��u��Ѭ���>���tW{�u�;���\ON����=lO&:�`����{�"y���þ��UM�x�� �6���_k�U�zTw9��)����x\���U���*�Q�Do��~jL�Fϼ�Fr����R�y�WT��klLbB6e,�v}�Vx�4���sR��~e��8�fP3k��Kc2HZx<�CV�o�^$|��*y;Y�����4��y����r/u��F��N,���d�AO���M(�N�o��b!�n��Ob	W�8�S`ҹlt�k{��c�I�tCz9��v�1ـ;�*ɛ��G:$Mhoo��.2���\�ԅ���UI�|27�X ����v��wѤ<D".��[�Ҋ `�4�F��Z�Cx��	pU��\u#�p��w�{���|;&��Rf�jO���.c1z}guݕc�# ���0͓6n^	.������݌0^� ?��U4��Z!��M?V�`zhPf�ee1�.���RY�H:32�{:;��t�!*�(@��=��K�t���J�tv�`��y�+��:E=~0Spd�a���?CO���DB�JQ�z+��%�L�e~�Ҵ/Ws.��|���X�X%��ure���r�V��Z�m������&ki����&��#�`J���E���oZqI�%eGR~� J�V����q���}aۈ�_���hC�H�����Uf�U`Ō)0���`�[�ח�7N^+�R�ۨx�3�	Tw`�Д��~HG�~@�Ξ�n&�3�eVÙ(�����rJ��1���HM�f6t��I�C{	��|��´X�"�%܏���j�����'�*Jӳa*1��9��ZN���|1���y����8��Q�5AO.գ�_�g�o�I��s� N�.�,�!s��ʑ�M���5M��ZO1�Y�i��qs����hE���0GD���|V�si��>�aOe��X�.@<V����}!L@4�R	O�D���4�����+�ݒ���8��޸�Vծ7a3]�(����p\��P	8`��BD�!J��W��f!���I���e!Hۋ���6vR������s���"�ZѦ�K�W��c�����}�x�de�CO"����LJ%�P��U��Q2g@��J�^�Ō�4����m�iC3 ?������{�z���P��B����7Gu��v��\1�=Qx�0C` |�; ���Rm�3FO�;����M�EJ�|�/#4�"��nڽe�҈���O��笢=�e����xT~�A�>��Udxk�!�1�X�:�#�:
�)꼻�U�t{��2E��0��/��1@�K���RK����i4���1��&3�uW	�@;�_��xE$��:��~q\� [�B������}M_}]����.�E�{u�ALd3�l�W��<,�ӰO���ʦTY� M�&$�v)��L�X�t�z�]��mgo��^KH�)�Ч������r��	�2v��� N�;v�,��D��%B��@���&_Ϗ-���&�fT�)`�>j�T�B�@s���%)R��,a����rB�� ?��ś��� T�ۜ�YA�v,gwZ��d<1Q��.�/���K.�@M���95��m�q�Bh��Au��x D5��8�lѓ��奄_��!&����䴐f��0W%�4S6{	
���M����.��Cܙm�%�t��F��Q�o �#�ؓ��CU�о�|��K/�(9�݅��Kg�	s��+�Sys�=Ah�~���QCZd՝���G�v�e����'������آ�������p�b-ĕ��a�u�3/i�a�A��J�Ĺ`	̦t� p����ί�V��_����7�\��q��ѹ%�d��o�tWE|u64AG�����\��8�y�JV�M������qHj��.��Uǜ�<�/�9�E .k�?mu1��M��# �K�s�Կ�^U�T�I�o�|,Cs X�DKm�'G���"�m�ϰf�����}jj�
�Ԣ�<�B�^F7�4wC�i�8=hXbHz*}$��!���ݱI .�\s��5YO��������s�!����0�3W^>�R����K^`����)X���?�`L@#آ̡$�)��+�*�w�99��?�x>�,p�~'��M�0��Z4Pچ lQ\��W�rk,bTܾ:�XQ|��ݤ�+Ű�hBpU�r4����7oֹ��$ǭ�J����k�9��;��P�x��@����,*oũ6�ϴ3t��d�:��B�"8��G9yh��'�C��ř���qf�gM�����N��@} �c�3P�Q�"�<��P�t6.^���S�6������͊ ֊u�h=Cf [i0:���/�$�M��_�������@�G3�k���޸� �G���3�j�Q�L>a�A�r!�~��7�v�)Bo˹͏�]�f݉z5��aS_=�H�����T��J��|��J��m>|��o�i�^P�I��e?���o����ꕤC�K�Ri�]t�¦�Yc���ZJyw��lݗ��$W�X��.b����J�ޒ�a��ߊ(ު��l�iP�� K��lo��+�hmZ;���n�~�%蛒[F��;����*p2S�����.gƐK��9��Sځ����4Iv�1�.?���2Յ����=o������#��
$\�k,˘k>�A$�_��
G�V_F�Z����i�d(ANvvǩ�l�\���Y|D���_���f�Ackya�yC�]�sr��C�N��� �*z��2A�6ɡ�r�5�A�༟r�[;�K�����ⱃYia`�ce�786m���aO�r�u�P˱���!�nD�⑼�sA�ܙ�YYE�2��Hw,4�;�*�>�@��21��G��p�f:���3��?lșNK���]�r(hx��e�o�t�X=���
١^��Cv��>"�k5�����g�$;g:�Z�ngk9��T�=�AԐ~pc�[m�[6E)V���P'�?$��
�� ���?`��W~b��T�@�+�G+
d�'��Ù�_p��q��
�r+�����H3��!\98�|ې��=ɱ}�2dע=��{�V8N��K�EF��ү���T���wfb�SA�z ױa��5ɜ��7�:��M��b�w�{�7&s��Ug��&��4�}(�L��E�ȫd����A��� ��W\kK�l
3�~��[���g� �yB�t�w�=k%qh	q�s��S�<�ģuϘ61��HOJ�h�#@x��Ql�#�eD߱y�c�FV]-�	���#U}�J�Í����;G�X�U	下��5i9�Є��t,�9^I�0vp���G�h˯�S�vV���'����[8��h,�+类�ޑQ]�^��̎�*H0"�wJ9�	J��|������+#6����~�6����da��^��dWcy6��=�X��Cq���(B�#��H"��?嫪��G̱�nk�+P��jT3�������T�I�]Sp9�:e����(��)\%Y3Oፖ�oH�a��;YB0��H1 ��hջ��.U���)��R0�;#�@��fU�Σ�/uT�Ka!���?�N�W�^Q�U���g�		=�"�s:�D��.�QvH�|fB�yzY�k��`�Ɋ�,�-�`�8��x'�u]���l�;;�M�j�<��SP"����Fh)ra�k����6�^��G��6�$h�����6}�����Q�V�����vP�De*�e3���I�,=���RJ��bA֘�M�:����%�
n[��p��j�Q�ڭF�$+�f����,J�������cC�-��`�τQ������	m	.��O�l���֊E/{'R���IZ�06��D�#�b5����/Vb���N˱������k�T�$(��ÓG�@w��E~�	f�j/1�8�	M�m��\��G�B�#3�U�)F܇LV���*J2E��"#�k�)�����.m,1�E1q�k���fa�U�;��ETq�fc$��Yn}�����h�����Z��I�h>8���!�����r�l���gܑ���=�XHQ`~H���@���9���F�{��'��z���z������3�;ę�hB�޻�D��%��-&H��-�q~X��`����{�@s��+b�7�İ�Rks�L45&�:`��}�[�S��h�$��tr��E�M��+^�����+�~�y�\��m[k0B� �lIŵ<H��H�F�Ƀ�ķ1k�g������I,0��҈-||�5��|�.�;9��@ª�j��ȂLpځ)��Ù9ii5I��O�y�D;~D^��%�<^/Ck�{�58�
�R,wjl��Y��,���L�C1���^.R��!�����{?�˺��K!"Y>�\�ݨ�ՠ$��ꘪ���d�:%"8;�L�L�0=��a�a^�R��9ީ<|)Ԛ���g� ���W�$ql�]�v?��\�d��`ŜL�.���h+�o�ІΜP�:A��8��# j���c�׃��;}3�������؎ב�x�
�!x�d��<�_P�b��: %��Mh�������5���l���G�m�l�&21�m�`���hޤ�)2�O'vA�]�<B��V0���w\c���C�di��"��bR*�Czˀ������|�L�����v�ߥ�'܍���xcPM�Χ���:�^f���U4D�YB��I�Q��L�3��i+Ƹ�ۥ��ϯ���1�Z4�J�}��m�EҰ\kut������S��3���W[�t�����pL?bO�����{Uv衎a���Y�o��qyD�Ii��٪u��n�~�6m�� dV�S��&Z׎�.q�n0 ��Ȯ2�Wi}������,١�����U�������e'=�qn�� �.(^Vr�%���x�B�K��e�}��\�h�R�