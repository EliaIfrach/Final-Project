��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$RU��Y���Ϟ�5(O���<��M�M�*<��2�	P���吏���}�rk�E3��⫨6u�Ы����<��V��52��V���{>�[�@��J��/���'H(N��W~F��vF�e}>8\����Ɇ7k�d3t���)�I%M1�Ɵ0����d���Vw�:�w����<�?i�ok58g,
{�!_(�
cZQ*K�]gHGF�ь�+�IR�Ղ�,mL_~���7�����(��%@
Õ&pS7��q�G��!T©V���rE����G8 #�+�&�)PS��|ȍd�A%f�B�%���ﻤ�����8T#�nhH��#"�ҩgzwv8��S\L['NLC٭��v��5>#�P�|с���aH��]�_d���2�����d(̹�X�DT/{|�/v���<W��iLˠ�Z�wg��3�3n�T�0k��#@y�$�TP�DK��d���KX��>�9��$o(�%������ۯ�,[�L�I�V��Jܛ��mx� A{�
fuY��,�r,��n(m_1��u�v�Q�|Nd"P��v*T�������r�$��2:����&mA�y$cv�b@W�x<�P����Ʀ����^ڎ�LW��U���[�@���)g&P�n�=����`.8��	��#*��m6 �F7�%ɻ����޹��X_�7�At'�.�px�����=�#�}_�"�h��$��m ~��M�2-���|����^d�N;m����-.����@�IN
�W%��C
m�xf���J�������]g�3�")B��D���0�R�E�E��Rj ��j&�c|�Ov}��h���]?J�d���1lV��T��w���t<�ʛڅm�꠬�]ѳD]g|�]���P��c.5#�ZkjW��G�]Q������i�jE���0�
��J�
w䭺��\MLO
���⿅q�fD��+�m�M�/2��%	((�`�� � ӽؙ���b6�>���}T��tL���1>�,1X\�&fe�@G�LL5Q~�W��Ña�2�qѓ��,L�/�sE�z���I�)b� �0�a�G��Gz�A<�����zSIܙ�I��dCǥ�O��<�%��|ľQ��zΒ��H��	_ 7W�)х%�߱6ĥ.C�Hr�8q��	+�	x�|e��߉���?ܘ�L��n䵭���̣���83����W���P�j����4�W�^T`�u��l/�պ�ӻ;��j�y�gP�F�t��ǝ��ك���GP��H�.\ �[J�bJ˄����rs�����������Ŕ��m�vťRS�ܿ�*ĺ������s�������cgi���N�ȥ����/?У��1�OO���R��"h_-����x���(��T"P�ݟ l�"��M,���ٜ��A���ˢ�M��u��0�=K�X
Xr�ڴ�QV�R�d��88H'a�]�u���v/u��Dv���@��:Q�v�����'C;/�nJ_����g>���WuK��t������?���P��c"*���޷^>19(�T]�VYw�c�)���D�
0vJȓ)Ofg˺�j9ҡQ��9ѝ��r.������Ǵ��6���3�}����9þuӵ�2a�Kw_#yI���C��p�L~�E2JŴK8��Ɵ#�.}$:�P��ͦ�b0|����U�y(z������_vp&ɭ���GI��{+Ǒ~�Si+�1x�|�
��	.*+=�^ef�!}{X�	�I�/�7����������"��f�L��������eL!<3P����Y:��Fv�~�2dM���P�����<��h!�*캆M;�
v�� �s��qS�ӁW���\�<E@�4[��-�(�I2]��p>+��Z�O\Y�v+�n������U��dd� ��i�-]1�Ӥito9�)�����&;,�V�R;��51#�,U,6@�x��4z�x�fO�Q��w8�/p=�F�Qc�&6�VM�s�E!t):�e�V6s�'{ء���l��N����O|�e����$F���OT�}A���2Z@@�ɬ�F��x�J�u"��W!�u�{<|\��I����8���c�C�}�S�R� M�J�ʈ�5�D�$��ȡE���������m1�!r�1�7�zĮ8.��"H�M0��"+E�	��(��կ?��R�jg���4I�.�C�?��j:V��Ҿ��H:�9Y����.�w^5젶�[��<+���	���j�2�9��u�G�*"��8�������V�]�@y���@�0�ɥN�e�KY)����_&%��r�A(���zV���Ɨ�����������3�,������E�a]R�������-D�D�ݖ�β�)#(?3V����GZ~ 
���%u�H��ۄZ8@3�O8TEX����cD��s�p�J�zn.�D�'��Ah6�K��m�T^e��+?wS��,l�TR#�&4�J�t���ރ�����C�����Y���ař�H���e
��B�וH�;>=��^�{>������O����ޖ�_:�	Z�������g����_ih�Y}�i����ڡ��3�75WO&�_/\�0���������d�ȴ,�u/�6B9��X�q���kAW�7c�W?�VJ���M}A8>;m������$vp��c�M��]��햝��+��Q��׬
��IVo`z���ԃWE 0F)��֢�Q́�א�QN�Lf,h���j�hÜ��U�{�Q�׽v��1+���D�,���
���Z��4��*����Q�����H�'gKߨ���t���"�۠[m�^i�Pl-mv��iN�D��G1�i�H������G4K���-�S�b=��[C��प־�;�/�6�"���3Xض���X�ao�y����<I��:/ڻX�*=`T����Kj��9����8�E�gqcp:�'�O�B���8����ֈt�cGH��,�EL���0��-�����1؃����>g����<�А��F��j�;L)�����WN@�$�>:��Gj���a��1��O4w]��ւ;ZB�x�S��*��m����7�_g{[]kڨ��GD�V)������o�ҳK�C.��0��ǜ�u�B��X�K���o��+=��s@�Y��ܻәt>�w6Wag�o/󋀨���p�=k�)��]��k^x3�X��N��[4P�V�Z0��]���Qͯ9=�_Q���s/(Q�E���ID��Q6�튾�Y�>��oz�J����z�e�i	��l�R�ȋv
�U�]!��*;��T@$b�bz�PlQ���-!��]sMd7[�����7���r�&�K�_��UA�C/|���n� �����������^���0���	~��Å��P>�3��|��z�aKݕ�z�u�c�XdY����T��oԿ���������a5AP;�B�+�%=F�e|0ԕ���=x�;D�f3�4i
�)�n��:����B4��V�&�Ct=����Fp\�������	�˂���?k���]aZ��Q�������ӽ�����8Z{�G���ؼ�B�*����U�y�	E𩶿�M#�&|}�D	'\-���HT�!l; z~=o�|���i�����7���Jb��eS�Ԓk�m��F*FJ�c@�18�Y~]��<e!r`�>��NIZ_���ho���^�þI	n�~޹Af�%@�U�j�jK�*����TA7¯��_#���Y2I�})!�r��6�
�,ƾu�p�+v�E��L�$����smI�Q�6)�i�
�ث�RE�[I�$�vΙ��K}��0b��'�K��P	�^�h�!vZ*UW,~���2v�}g(픜���������<��Dh�u���'�QT��|.l8*�G��5�v�q�cOcydZYor�,z��c�-��?u|��F���-k�Pkz�)@ۂ�EI������<��a����b��,t¸�94�d�c�L_�l����Z
�2��%�����yhP�b��[\ck�vc�3�PQh���k"�x
��>�H)D�!K�6��-|:z���qA�2 �CZ��#n���+��
9�[�_{]��`F3+��M7w�7��۠���e�㈔�H3�46aTz�ȏ�Z�mEɬn>��BVH�0
�^wB�-����d�&�d
��07��;��g}���該����=n�&����@p[9�ի5�q��q�[�H�鴣zK�i5�R*�p��8&"`s7������D`�T��itX�J�g_rJ?n�3�y*;~�.�<��)�����I;:��7���Qr�'�R�����dxY��H�b���z�^uP�;�gQW�=�l�Q,���4R��/���^�ef�����C���05-u��N?OZP:�����in�W��!Ƒ�px�Dlb�m�*��	b�Q	�c&b�!���O�C� }�N��	�.�g��}�b��&"� ����<Cl�J��^K�\���ـ�!�y/�Yr��8��5��Tl�~��ZϜ����2��N^e����x�	��O.t{B8I�wT�nQ��5�#𓖙B��8P�c�(dfʒ�/_M��K����K�i>��nW|���n�:-P��ɹ���T�}��L����hO���m$G�k<�>df��ˁ�:x�B��J�@���9�UgY��G��Q%HkNo����&uTk�<ǒh#�7�kjMAPܞ��̌�8{�T��W@�JC�`� ��W�(|F[�Pg9\�&M����aC� T|�?�r8C�{����1Q��fc���K�zt�M�h8�}��B6Q2�߶� �W�%EZ����F�P�y���'∿�,����5>�&�+<o�����4�Ґ�d�^���������d���{�W����.��Ǩ�~�#�*10��JG�)e����D���[{���ء��|YJ�uʫ�W	ö��&�~�*��b�u�)nG�tW3��YS$��-v��/S(7�՗q;W+b%`b�o�	"dB��;���řv�e�(��ޗ�qՔ��U,��s�m�d��᷎<���r�BZ
�.��o_ߝ �H���M��[V������S�Z�v2_����,��i�<Е��HI�CC藥��܎a`�O��W^� ށ��N�ꒌ����Z�6�G����)MJ���� |6֌^_#I��*G$�D�|lM�'��ۧ�+�����/��1�)`��/yPwj���.s��
��OGǋ�瞺���7�.�S��w7^6Y��LH�>���5=��u J����<�4г����E�Kpl�������+��V�����~������J��>�e�9�r��Q�c\�և���m?a����<��f{vUItJxr����+��*�"f����i�)�u����3�3E�dߓ���8�"^��mZ����eB�́���ͣ�mXS3���,-ͦ ꍖ����ƴ
�I.m�=:G���U����G��S����#�q=�⑐�A��ڼ�LY�y������'ױ"oa��M>򞋴���("����Ҍ؆f��c�'�rj+^I'����t�Çc�d��P��;z��q��&q\�1�,�^����3��/ޚ��s���̑B��������Ll�
��ǎR2Lxj�U��X��e76X���+N[�A<�qa����,8�l���D��0��3� ʚz�Jt��H�te�@��L1T�H�l�鏯M��YjX��'H�	��w@ˍyR8��Q�-�Lm|4�'(��#K"d�ǵٯ���(�N�:s��ۯ��(��`tj(�`� N�'�_��H�����ѡP���b�s�9'I�E����1����c]R�4��`�xj�w��	|�q�L!v�D����R1!=�n�L{���b͑Lp�}?YM6G���N�뱾�[��+�")���u|�c�]�ܷD+^�iI�;���S���6�����C�0��d�Wa�O3VK��)���X�D�D&���o��M����f��Ō����Z�賄(��l�/|4�)��Ʋ�� �N9�,=Yj8�v�g��6�q~
މ:~�B: RzE�����A������na!�Q?��̱-4��=�&���	0�Η�S`�Xg�u|�[��� ���Y�������o�OzU
^Gf�5K"xTs����C�Ec��9��IԆ��D�كBM�/����|�25%T&w:�W8/~Ƅ,�uv��0��c�&s���М�}ǁ*Ptqi�5|U������F�i����t�?K�)���R�t�@�C}R�<f�m2�`�V�ƕ������ky��%�>���<E��b�4�o���nC&�N�$ńH�"0jj��'���"��k��?a�5O��M��Z�ܜ��E��	x�7�R��4����b�YʦC����j�L�j�B�ă�k2�mA�$]�l�(��%�7��Uȑ��Vn��{�cg<	3Y/�O��#<��=���_q�Z\�H�9�wO�ggL�̹nܧ����h�V��=*��2�>d�|��`2���Ǡ���j5�E�H��(�-E�^��m��nmՕid��1����O]�~i�#�i���RdۻBR�j���꘰!x������p�DE�3`�_�^<���������[���a��̬!�*ۂ��W���͔�Ť���h�o5��4�I@�b�E���D�5�b���|�L*B=��X�̪�-�6�D�n��JDμ�ƙ��������4��3&�6e�o+��{�a:�B�t���+�RnTa�E}����Y��NU'�&��RBt��Ŀ�����r�y����P�8B�jǰ}1��z�o*���:��e�����RV�~�-�+la2hЛ(G�����?�(2ۉb���!��`5��dWK1�rG@m!�E82�����YC�l�Rn���X�3��g��}�o�+�l��K���]�O���uY�f�9�vPH���h`�}����hN��Ud��_��w�f���q��1
10�����r�Z>w?��:/�����p=aQ�L��o2�jDlfb��>3f�$1��T�A6�"$U�����d�:A��t�X�ezA�@+��h�2��hYM��Sx�F��I��B;疪ad<��l�����S��RM�� �/P��JYȤ3�B�L�s-�5�����L�v��	���@�[�$t$�y��%����5�'�[kX�4/�l��+�s�[���#�ҹ��F��g�C(8Ru��+���r���.Ԥ�>����-����q��N~\��R��`*oѬ� \��N1�o'��j��KC��e�N����*Ȥ�4X�|���*ٹ�vg�pй��>3Ŝ�ʹ,���4O�l��R����P�S��ei�E	uO����'	��"'A}m&M'�]�JI�L��p����^��wWuHY{����+;����k�b��2�E�V�sA�gc���\
D�D�Q֢�9�4�Ф��Η�(*g����㎎��r�n7+X8-{�[��a��<��\)wC�"Ì�{�-��,k��?�L_֛�jT������f�Fۓ��e�`�!vId�C�<$��m�V��9r&�M��~5Ux���B8Ce{ �l$��K�`�c`L֫��Τ��O7*.B���͢�K����ȓ]�k��>Y�xOSS˿�!���p�,Rk��3�/��lv�X��W,`r���όt���ɍP��5�d�epS����%>�"�ӧ���4�����F��Ц��[�bFxQ�#,x���r>��\a�e8�Y0M�TO�;�X���3D�lA�����0�\�a��;��.���n��S�
;�x�*�f��qR�HŘ��3fi�P��b�Ͱ�}���g�d3�sW���[��~������{�:C���!}�]���b|�?1�mpq��������gm1�&�V�|?X�j�X���p�8�P%��R8���"���T`+���|���N+�l�����MP,�Z��;#=�&w��&S��$�v��c��*9����m�����y`KGN}Msf��:u�N&�i�Ǩ���D����K���_�u�'����h�~�Fɶ	�M]R"�b���O�	�Q����t&W3�ӹ�����כT�)q�hc	U��Of�;�;c��	�w�Y�oj����%U��0+�t$T�����Y��2�H|j>�����ďX����!�����{ɲ���	�z�A�si%<�($>~J�ws8"_�?��o���A���VS�I��'9��kĶ1��t�6����)0����~�Z�|�P���/a��Y�U�ڧ�*���҂��hgX�#j��vuZ��˶p�<�"{�PZL�(�6�B 赥��P�{�l����R��0��`?�d�r��S���K�ֶ#�usI�tJf��ШXi�U�M-��]�TT3�S���L���x(��uIrt�2�Js�8�W�n���a%��" �2�qj#���P���tg��啴`,�#oŀA�͆��o��w�V؏�����l���8:���5K4��/�8����WW����R�n��i��';����&�z����>��y⥉�������-�i���\��0�3�9/Z�".���
Ck#�-	3��b-_�5]�s�e�wi�ϴ�O�*  ����ź �� a��  Z�|�<�_�z�5D�����dG�4e�Ƅb���ݏ<PW;��׹I5����1z{hL��0�_2��W��I�/8|��u9|�h�)m�W�򀨍�i>|���'��J��ӷ�\�ۆ�؁������NY>�Y�!��D!-?j#��a�j{o�$Gd��Aw���5?g��L�MW@#4��S����r�I���[��]��.-`�V�����k��ފC�rb(5��'�����R�-!y�E hMj3m��1ނ;�xY�`.�n�v����`���=��^�\Y�T�`5�9�S3�������$wiA�)\��ƨ����V.7O�������ާ��ڴ.Q�����߶&��q�טJF䯳k��K'!w�[��C������2��ȫ�!��4m��ka�r}̉)ٔH�譏��d���~�0��8r�Ar��+����3�&���q��T@Us=�R����(�&�!X&s��8��~GcR$�X�aQ������^� ��|;;�K�WsQ���7����9�D����J(�7����*U�)���/�4�"J8���/{�w�d���#�1T��ĉ7�#{���s�:�;�%�(�O� �۪lо2�:#�q-���lY]���-p��j�=6����-��z|	�C=v�(�D��9Q/ة�ł��l��v�&K\��SrO�o~̪�Uf�o���[�xa:kF��cb���*ⓗ����4冑H�d�AK�e8Z�\�9uQcrݶ1"��p��9g��^5�6��h!j8�2���L{��J��	fc�'=|U�w�#�SM����-1��ѩ��}!l�~Y'At>]C��X�꤉��덾2�!*�	�[k�U�+*v{'4�;�c�Cy�QNf�Ƈ�E����ĥ�~��b�U྆��o'.�[6y,S�RωsY�K�K6� B�T��7
�8_�:@ܢ��aTf.�#�C�t�)�JӽH�����s����;E<QO	��N�,����)�ܹ���T�����-��#��x�C_���Z��a��/͢���Sf�SH'-X5���+7�~�޾�mβ{�����IR�T콈�_�ፉ/"��$R�qȀʈ�2<z�H Q����WI4e}�76��zϿ���&!w��.�*�� �=�<_�;��W�.yô=�J����z�8��e�;[�:!��z*�q�7Tz���S�.8���$�G ��֒�M1��ea�@M�C �8�c�Z�c����ٯ��d�nq�����^��y ��K�?�������F��:���N�lA�_��-�jlBvd�%�j)�#H��T
��{<:A~r�E�|��`��𕢈R�H_H3?��6�}����&����f�LR~�W3�*l}�KgN;$�欻�9݅���!��#���GM�A:o���>���3Y6�r?NNu��R�J\iv�j�׍Q��������CX&�c��tzY���нo�A��SĐ�卞KFPd���{�� AE��A�����'`b�j~���R�����=�v��M��k�+�y�,n`��`Ƕ�B~�vL9��xK0�N��O(8zkl}8>̤Yze��{����3h��^���q�N�� �5k�[�W�&X���U�y^�8G�҈bwݱ�VR�0�+�z��N��9�(U�	�V�զX��T���7�b�A*;g��נʠ�nn����*f��X#mȄ}5E�Y(:��3ZvC��7�%9�ڸ�a�r��x
e��8��#܎M�m5��O���RG�O ���wa����%��� ���$Ю���M�Q��ƅ���v�IW���nY�<�~�/s�"Ő�u�@^#[�̋T�Kƾ�U`lΌ�nؔ�Z�7��G��:�?|�)��%��>8�5&�&K45��ߐ���E�n2��%\�
G\ U�
U�%���*�C#��vv�Ǉ2�4�ģ���6�Ni�)j��0�?��;t���4�x{%���.S]?���uUl�����OD����!�ޣ�����ZYz�j�y�S��� KԴ;	�ڀ'1��'��$�7��Q̠�H�ʆ���c��ԡ�❵(RR����v�����~X{��JJ�D&$�ݪM;&_\6�1?_����f�wBA=D�|�n-�C�X�Pu��UDfBs��v	�$'D��Uj-"h�j��y��:p��q��i�{zK��Ι��)E�?�$�V�B���Z7�w��t9
!��[�Re*�;��B���~���}(��9eSw�LG���|�_�K6X�����$��I�a�&���MI�~"b��O�ܴ���R���\�8D	�셗xq.��_���N��L#'���έ`��@�(��plP��M�S��׉�*����i�j��Āi_�)侏�g�RkN��3:���INtK����9�M�\p1K���.���Z���fA�Pf9���+p�`'�����ރy�v����`�t����SBm��'��f����I���-�.��J�]�Z��8%��J�>^���&��w�^i�ZUk�#5��L��d���/VqI9o�O�*�>ʣ�u�	>��Dn�����=hub����*|1w$�x�����T6�ď�Ddjl�s��:�a�Q�W%�����u�ܳ`E�b*I1��_rL�z�C���t�,Ԥ z2b1hQ��H-�F��髹�*�誼M
]�[ �)M�B���a-�/{$ϬDV�w����3�֑��w��zŁ�W����:���2-�YJ	A�9�P�ew6L!��r	N�Ű�#0� ��s�Z?䇱�� ]��`����q��Z����Z��*�K���&gR�ϸ�d�A.�\N$�T�Bo0�5�� ��~7&v5��{2ek��}�br{��
��S�5�),�q�4�W��R��ײT	����WN���Me �=N�a��}=�'��Ąx�ة��n�5�@%��h�g�~i��
�����)0��9\yf��+�������mwێ̬�5�GŰ{X�8�:�W�2!EW���}�A��(g�{O�,��x�7,�P�#��$t$�R̿��b΢�l�l�[Q41ݍj{��<>8���+���t}�z�X�����5����%��4�\N�FY��N�Y�b��z+!�6�%c[�����iCC(���/ƖeT����3�,��>P��3�|%>O�M�-�ҧ��혆�����Y�DDx
�%�[�����؁���?[�w�K�}�CN��Oѳ�&�g��X��ުN��T/�ȏ�8�$ $�U��ZIa��2q|��:��{����l���g ������I��8�����
;8F0��Wz���� �i�P<k|�4�ƥ9ʃД��%<H`���rp'�%}�;��9n ٘ZQ�7i��Pd��q�'����GL?��
�/햒�G�������#hۓ��c��Cś3Po��c�o=^��y�T|��
�O��Z�Z1���ci8���L��>6��)64��qEe��c*��Կ"(�ԵQ����% Y���'��s��G�R���PHİ��O���8Xr��0�9�U
��c�9*Ca@���Q�A��J2���#�����w̷��J���ު0xBUɷ%c������9a���ͳ����+p,������V,}\�J����5����}� g��0�-(�7����^��H��Q]u�]�Qg���i�� Ae�~�_@N��7�a��ӊrP0��n�	}��_���6X۬����lѽ(�m��&���_�h���'M�W�ȼ:T�[	n�.v��`҈q�F��d�l1���:!l�����6�6��՘�4���e���������u(qǨ�Y�E���)��Nu:�c[*��H��H�<N�!J�_���b��g�*(���@"�� ŌƵmG��Hn��&�v(���b(������);u���:׈��z̮IxO�~�ףA�AB���ΌΌh#�	ӟʩp�Ou���@����XR�s+f��0p���ɎS�)�S�A%#�W��n;���>��9֣��,~���J��6P J�f���M_l��y1OI�1��Th�]3	�.�=y)N��M�M���өg��=M�z�%5\������[t���y@���������A+n��c���+�掬�Q���4����jF���ϛ6�4(ه� V�#���}eSgѽ��Voڷ��I��������Bu�Df1��,S��p���(�|&�p'�>�c���[W����su�Q�Rw�� ��dG�]�Ԝ'y�=%~�,�:��=f��-9(i�K�
6��A:��A*���n�ui��ÛI>"��S�Rdd���n�� �q1A��t�q֐���#T���k��	Ґ�N[pq_�k���v�yCǓ�� �8��Q7��-47�n�)hݴ����\��Y.I`�K[��"U_ϧ�g�KO4��1Q�<>�k�@e��P���?���R�� y^�'�ȥc�G%Q+��U(~��@>�v�n�Ģ��k�Ս _�o�{A��U�wu\C��X�u���{Kz.�6L������@�}%Q��(rQ���ֱ,O�N�3��t�}K;�%�=wH]Sȡk��|�G�H7)-{a�򙼱�c�}N��~gB���*|���YB="���N��e�f�5FFl�˽��9�1��<z�[�b`���>�0�I<���o��[��J���!�G��6|}��w(�7��b/�"�~P,��P�R��;fwJf�}�~��V`�'���7�	�7~d�`7�|T��GanI���X~�=^4�A-��u"�GE���P�Ty7��P)��@^��'��_����7�}d�2��d(#(� >5@��>���~��A�y����(��՝}�yJrі"�(n�\afX4;Y �ZDY�����ó���J1�UKo�g��$���.kȹ=��TeV\�;������W�3$D�q#d��-�]�lk'�������A/���g͙�@G�:��q�YA��N��خ�MadFd�{^ϣʿ����t<ħ��;B���+����{3��	�{�֧bj�=���<�Ko��~W���p�p��$r���m���5�#���Z�T���|4�;ࠒ�t,�n����Y�Z��#}�Gk��m�� :F��d�"�*D�zQ�� P$�Mp�8�A�T�y���ܚoz����g/1�feC&67���R(B��#�2�I���^'���9�hn7'�a�_�5Ly-m�H�$2�6�r�U�����=�9kHv#�+"����J~��R�m*�1���ebw̚�kuOOq��-@DE;���e^����������r;�ډ��i�Ϧ��v��q�ShP\9اwd(���tFYU�C��Za���]~~6V��}}���l��WW�:���A�L%�5_e=�F�����y�p�ޯ^���ƇK����6|�3*E$g�]�����#��L�>�$�����͐>.Hx��@T�+Tn��%r��E���f�4����DE��oCE/������c|�������7}�4�,�W��뾒S&?]j�Ba��N$m���
@l��5O0u!X@��,�n�*��+_X̜剾��m:��G|LL�D#걫Մ����1���fu����浤t��U��3����vw6��,h)�f8r&�::�s+�14�ڙl7����L0g��=�~��wn�TvS�0�n��U�瑣����0!o��4-h-�n+��OB���zy�)� i^hX�0�m�	��٢L�V����A0�����GG|��j�t۸iw7)Z��M�>$�h��\�>�z�=�_t�X	����'�(^����œ�ϔ����i��XҬԢ�Jq��0655��m�{����� ���Ն �na4�袿�3��}A���nW,�������l9������X^��@&R?�IH:���P!��+�F��05����<��ɦ�aE��@l$��n4�v�ҥ́J�.�Gk�xN�I�{@���<,�b�PYǒ�Q� ^�j� ۣء��hVT:�|
#�
f�׷}<��ߐ4�\M�R4�▝k�U�%��il,��=9��x��ķ:=k����J�O\��Z�|��<�]*ӳ��1@�����'N%�O�9�EJ����`�����8���e�� ��5�Ҭ�N�AG͙���K�>��J��,β�u�b$�m��g!�d�h����<kdO����id�W�3�5����J�SE��3��^3ޚi�,�\38��x�4��w��_��UѳV�ޛ�UeZ����ڋ/b�Ef�k�L��>��DM�F�[ng�	����#M�����9�]�~�s���;d�;S`����o��u���������,� ��9�^��hQ�Ԯn��u��>���g0
Q�js�<�b��"R~xm���fw��eFB�?"����n�K8��8S$��i��4d�����ɉ�T#2����K0�2�$�Ž@�����.��DFW�hIw���)���Ź��n���f�t��a�v޽��.�g̴�����㓁����jR�`�DX��$F��4e���#$�qU�rwxda�s�_�jg�	O;�0!P��[�Β���Y .R��hQ�O�S�M�0�&4�/`V%��%�.��N+f����izi3�v�a�p�*\/@�{�B.�,g�P����nW>��Id�Y@�_�RG>�s}ӽ��5��XE�wF�!�1�(�=w�߹���9!�����+���@S(O�@2)�F��h�Ѩ}8�F	�Y��1���ґ!�}�sHa�nw�<�a��U+���7�`�e�N3E�a;oE��2b�B�/rn��q���WJ��/Pzf'{���oj��߁�(�N������3Z���ց��A) �
���}��@ܬ�r9�U��`JԱI���G�w2�񅪦��r���������¬��}y���:4���Y�.��ڠ5��cvЫ���e�y���[�Bv��ݍ�]&���;�̪� ^Aj�V�g�7� I���x���0\�G��$����%;�<ɣ0K���(Cߣ���v��~�ݭ�F���\���������cҠ��qb"`�	��:�z]�y�:��5"]��At�H��}R		�D�`$��U�oP�E���@Q|�l|}Eg�-&��̲��
r�r~qՒ�YYA�V��a���-⒬�Z�ҨP9����̕�Z�����0�7]��p߫���\��͒F<����EYp��d��tB&�v��,O�E�y/ä2���SK��=a��9�� ��|�۵��js�7�j-)m�Z�-ɣ�*eGEЎQzw�)l��E�N� a.���s�k8@N�b�{^{Ч�P�׸'y>�����B�F�s��H�`�x<5��G��U���ky_��\@��9br�J���1��P���Y,z�4�_�&-D���R��HY+�O���*�K>M�/Җn�
Y���Թ�z]C�s2�jm8o�=PV������k�o*AY��*�
SX���w��Y��$��P���{��{͂G'�$�~�K��S+��B�έ���0�����S�Dw4����`�JU�� ���q�����zm�J:�+�u����^��̬�4#�)��5�w��b�3c��_��
v��Q��'Q�h������}���0c71�Ega��RD���R�{m�{\�P��WA��f���fx*��t��f� ��~���V)��!���ޕ�/��C|K���VeՎ���%�K�?�3-?�3�|\����������>��S!?��WRC��׮X�`��@U���S��|<&��=X=i��!�Q�,�i��Rq���o3� +�L���qv�'��\*(+8�,{� K]�H�-N�6���V2���
F,�9HR�F���t�$�C.�9���`�QѺ�E�S!���W|6z�!�����Qοv���(z-S��|U�0�d�����5�3�Vȟ�f5C��k�7崠J>��J"�����SQ,�m��o2vkĦ+���� ���+��맮�D���G����A�/ب")}��Ŋ��}�A\kv��-��)^��w=`Ku��o}�4�xF�p�.����}�6�H6���~��$����2^��&�V�s�f�_�BM������G�(�ܑ;Wo�_ ��p ɷ̈���0�߈6Rmnm`pe�D�W�q�g�^<��n��|)�ٝɓl�ˬJ�v��c��O`^G?�o����*����nWi���{F�-� ���HoS�iJ��&Bί��-\t���J����׹׻��F�����4w�/�	��ݬi�-����"�G��֐�4��CEo,4�"��D��k����m��T���*g{�� e>%՞wDY�T�'��oԈ���G;[�t�n����n�ii\�'揦�B*O��0�:i�7)^�m�(�����~�v�r},4Â�,l�b�*�(y��
��t0֎�?LI;��u<p���ܟ��y�5�z�;A=����qۼ\�1S�����G�2?�-�ʾr{;T.��n���
N���6�љ��+4����`wݿ6�����V�]e��_��[��-�l�B25��+E_�S	܈c�8�!��(�3#���@W�y<Ju�Ѥ��� �7�ys�yόj�ul�<-��t@\w�wBl�*^��96,�l��<�1��������˧�S��c���~-��AC��v#�K,{����8�~
�T����X){j%<��ew7�F�Q4���Б��R��h���
��b�I���l�~?�h��*eȍ�4ꌃ���D�Sg��!v�W��l��1Z�B�g7� Y�FD� ~�r?�&�$oG���.>!Ԑ�!&���_Ő/[e��ש�'>���f�T/G���/��B6c�(A���� Y��=��h�G<ݵb�i<m2͢���5�8r͒�lſ������L�I|B=�#sܸ%��-|C)��#i�Txf2}"�剅X�ڻ8�<�vٴq9l��r���v��a��;~��z�>[n�Et�H�/x��>0�M}���4�wK�p��[�����
� g嗁�Tq|�N�+�E��-���J?sl7��\�w�1��w���u5�`�5������!_��{�Ta��:(��� �*Z���J�g�r�㚖k�����.�n�W:]ғߩ.�r7���`}7���I����u��y��97�+����<�G�!G���������X\`�/�4c;C1"��)j�>(5~8� �K�J��=׳����T���%�eW��jZ�p"iu�2ӈU8�;�-Ζ���iw��%�g�3fqca#L�u�h'��A�I�*�r� h5zjj��}�*R���]`_T8f^�63������G�L���Qb��N��1��{#~�g�#6����"&��Wc����g>O�O�al�I�M��^xu 
�������N�����T�"n�~?B���uy2Z>ݟ���_�cu��~JՋ*U��첮̡aю�!,D)m_��er�;��JO+1�����gH_�r�2�*�f�8���`>����M`�6���p���e+y�]O�_ȯW��%D�+�asG�՜�
�2�^oq,(W;�P�,���X����r�%����3�ɮl@�q�Ih{�x�/�:H�U��@r�A�Ih��HU�u0��~�It_����?N���9r���4j_������->d[�cx�H$�)��p]e�(z��߯�XA��T�>��%��R�VS�W��-��FX�1�	�:IĐ��D@46o�v��wWT��֘V$ޱ`.�6;�L� �O7��x�W�xT����x�"�[�������X5ɘ�61T����4wsv�d���M
�v���L̞ķ�χ�#��M)��i�W���
�kQ����b��e�MU�-��A�\b��0b�b�|7$x'��Fb(`E�I�v+Z}�`����J
��<�Õ>X>ysB�D��b� �O�W����&��,�|���Jeo���D9g6'��%�A�����'���h\pA�V�r�Ѽ����`:�����!���YI����P,��ЏN��s�Gý��*v��9���@�@���/��[w��� L��$��(.'��c.��F�
��"��䊷i��A�#,�p��d7����Xt��HĠ�*��>��{:I�Mȁ -!��9�EC�Sk~��~y�tFpRD��m��\d��C�_�� ��w��]�����W�"�o?9�3��N�P눿�%j��I]����=�߶�ٳ.�؆X\�FAȹ>���g�\ʿ0�1հR%�����PL�y(���(eB=<1��)Оo-��Ǔ-�M�F+�����'���l�T����K�=ɎW�-7��2/%�݁O w�~w�52��������.ӔF��ؽC;f�ocO�q��+~4�L,H��M:�N3.��3m�,��^�a��Qmn7�Y�q �4nL�f�۵MY�W�VW�4Τm���wIr��������N�-�~�iP�"3c��v�"��/f�&�CH�|T7���z*���6"s�i�����W
U�v`Wˏ��_���o, �Z]�"M����������q��ȑY�<B����}�i��,̍�}p��c�z|��ᆤ�<10H`՘��"I�R�tzE�4 ���>����Ո�;�������M�Y��� ^�Ȉ�"�&��@�?�؎�9��`��F!~� οj�wTu�ͩ�k�QM쏧c�BWo���h���2Xk��8�Q������C�4x@7`��*���5��?h&�t����լ%��\B��,Rw9�?��W��SV��V�>�������k���9�;d�*�U�⟟�lI�����D�6�T���`�+��O,��Xx6c�6_��v�E򇭌Qe-���*?wT�
=X�x
E�C��ҋ:ުo�B��*}�S'O$�H�[��|�<d�JE��!�����*	�gU��t�Hi1�8�U��M'��ۏЈ�p�ɳ�Nh���*=	Y)���!�:��U��I���q��{�B~��s=�ű�C.�G�轖�[�d��6�����.�jJ#~+�` ���3^�,���)��\������Q
t66Zk{�
��:Nͳ�6E������V�\�;�<iN�*\�>���ީo06��V�\;)�l�5E
����.׼�%�����C�S|�<<��ûm������!����O#.<�o����\�d�?����m�<n��tah�pv�����(l۞8�c�A���Rx��iy=R�өv���Y�̚K�i`�i�YB�A���r|&��|��p��fxR��Gg	YT�~��|��C�o�p@B���Y>$��a�1�����l�L��ca�.J3���R?��0��#�x����- �C�7���K[��t�s��E+���ٶ"ئ�-��(xL	��ũűo�g�;PRj)Wv�Mޑ7#����]��k��?�%��23%?q�Aз)Ef�1�N�Tf���ڏ!H{�lسmm�b�9�-reW)$�8w"��)���R���{��VP��
.kέB�8�x��T|�	�D���D��3�� �Q�}�.�z(�)NW\��UK�Rc�蝬��+���ꐊUk�@z���?2����|���c$���@A^K#f�Ѧ�W�}WD�yX>?��6�˞�x�ZN>�n5�؜(U&�U�Ů������`hti�	\cv&�m[E&�X�.u��� �ȅE%���0����+��e�@��4y�aZ�@j���t����7���t�N��Fӆ��R*ӦgyѪ��d����RO���@H�!k2�k�X}lt^ �W�"�X��m&/�2`���C�1I��1�����8��bV��MP��92(9
�����n=.U9�6�w��+���.5���릓����C
��{x��0e��[�-��<+Q�e�{"`�^q� x@Z����:��-�0*a7��m��U���&���������Tu�"�2����"������o4�^��Ȋ��K<�,��=�,�\��Ltpl�����
H� }�7rW	�εLp�������@v��	��b��B�o&���xZ0p��"�"�.�dS�$�h撇$>^v��Cӻʕ��=M���ԏ�y�#�HŔ+\cE��N��$C��T��x#��#�%M|�(��7��=s@HBI�Hv$;�)�ӡ�A��j��� 7�d6m��c���Z\���tf���� c:�٥Zӱ^n׺H�D�H�p�ٱ��`���sg[��]��� U<��ė��G.�v_	s���nNe�ǜ����m��Sp��R�J�2�1�(ǡj=�����x�8=�?�C�VO�+�DNOSx�qe��|���֊��/�6�����ny�q��#�r�����L���C�k�h?����کg��l��C� fu㤫r[K�+q��^}����A���懩��s� �ҡ�i��A�`ф-J�-�l��0X.L"W�2��~��� }	�)���Z�o�^�D���>����$h���}�MGֵ�ŏ]��|3m��D�pN'�O|{����l�!�c��"�:6����&�y�ڟ?�j�jr�TvMd�d�v��7B3�s)jQ�i����9zSE����:@9MD.���e	P�8��Y�R	�ϡ�ƚ�}ho�=��vO�z�=0<�Щ�V�S���G�w�J\�'�Σ�|x P��&��#FwfӸ��"9
�g�|4tCD�� ���+>~�������qVW��C�o޺�ol6�ac]�u���j��&�<���t��^M�S�C#���^���e�	��G�T��h`�
���.Yj>�e���T_2����=-�@�Qi��9� �m�VP�T�TOZpˮ�f�h�� ,��P1�
�~�e�K)�z�+A���b�/���dz�L���*A9�0t��'��t�d,$�=�c���O}��.S^!�$9�Q�l���1�=s��T.��N��E��v\����;n��?�NM\]����@��.�4�>�x�ls���;���Sg�f�c�A���;�3�	���DRʂ���1�X[������b�1i�`�h	�k�>� eq�'r��æ��$ȅ�� ~�o}Ns;�7�G����y}�S�����-]�T佚C�lH�+85��V�r�I����= fU=�ĕ�� v���D�Na���(�z$\��jaO?���� ��5�â�A���a.�L�K(�S��1$�Ƹ�&���dў^u�̈́�]%�R∷��#���X���v�^aYb?�Q+�`���p�t�΂��_[�ݼڝ� �J	�ؒ�:�`�K�l�
�؟�izx�q�y}��`T+�{�8S����pbځ��O-}lxe�C��d�^�E����>$��0��$�=��1��q��F�w��K����!�k�B1�^�kPx�,m9��G�L��|�f�F���(�^Ot��zD7Z�J?��[��(y"�����s�@m�׎0�P�ѕ������h����Y�!�! :j#�Hl=!s?߸;�rC䣹�h��8	g��I��ikE=�E�UD=E��W"�Wt�[XuV��F�[���+�#
���o�T��^�N�L��@]nu�gt��l�b������w=�zK��	����!a��:��B�t��g(K�l|���d��Q(�W��!�U�H�U��<��F��K����x2���Ȕ�����܈��<�%�&��9�P�������	�l����MƋ�� �eX�t�ֆ%fni���Ŋ!JV�����Қ�c�A�R����,EFpf
�+[-����w���WB�ڴ82�k�$挂�J�n�8�r�@H��u����7I���r�ou�$}n���^P�Gt?X�L�+�U�;��������EpT˃ɂ`+t�Hm��D��k�1���`��5�-w���|�=����.�ܫ�h.��p&��W����ԣ�s��o���w<I��U���"p-@�ϗkmn7t�-�eW)"�/c��?P�f��^���E��&��� ����0�j�P���V��Kav]����"
\�5Ϊ�s�P������|�=sgT��ݛ�:Kk�A΀#MBoځ@�I��ξ��(��ZE4�P�g
� uP�s�󵣆��Q�$��	w �i�Pr�Ш�)�P����%���{�9!�@�`�%މ�x���aNR�Q��1Z�Nv�[j�`�ߍI���!�@_�A��K���Z�D���n^�֪�;�i��3�L5*��W%wӼ:�
*�1H��h��k��������KW�5����Y1��ϥ9q�/6��:�)f��I0y�L�EK#-:%ׯ߉�
� l�_N��F��'@���xk���JSZ䜷�� �rb�0`HP~{#Ӈ� ��̡�IS���C�q�����H���/;��S�������7�x�U�,b�bP�B�)4�=��d�I����]����ա�� �0��4	�m[�W�[E�6�v'�1�(p,�M���(	�-1紣��?O�ћjg:��16�k5UƠ�>����ᩛ�3k�^���5������{��~�����n?��� � �$2�+�Ք}a�4�b�A�g�U�)��>?�L��u��!OZ��(�
{�N�**��H���V��s[�3���7�qX��_�$4�F�vBP~��W�n�5H����Qe�^O�8䳶�,�LȘ�˘3��um��$�Q4x3b��􏜦�c�B�H;r��K���#�Ft�r�I����{� {��ɺ�U��K�@��6']�VU`�����lQ���-/��cW��e?��U���or���W��?��<�4T./f�i���3O� �0���w��'��t�s��a[���C�x>*��W4l�����X��C3��̝~�V���'饱?�136G���K@ ��#��͸OJ�:����h��sY�����&4rI3�_�{Ã�ԠلYnek�@"��zSK_3nq��դ�Ssvm�~O��.�H���:��$�	�����](�P/BӊO����q�@R�ౡџ�~��~u��؇dS�g#�$��p�]�6�L���r*���:�G�?D.}��ZK�5�Ό&7;>Z��
΀a�K�^���c�!�,d�/4�Q���8L����"���;$],��뎓�A��%�1�x��I�ϛiQiz(�Nǎ����7�17�za���a�
���
�a�fL�Y�_�}�'�_�*ͯ&ˏY�?�K|s^`x�Ʃ�cy��Wq����,����o��JTm��"�H������T:�~�8�]I�A(Bȟ;ˀ������C �~�$����.+L�:ߏ��l=��������뵷������阳����SS��`�Q4%�e�
�v�}p�D�̝��'MD`1Ͳ
^
л6b��!{,�Q�{�}�}������&�y�U�@����F�7痗?�Ѓb�6Q2^cU-�z�I��i�����Z���S,��U��O�?I��2���:E��^�T.��}�(�H>t��&���u.�ɞC@W������(�y��C�B���(��0�T�[^³�F�.}ߖ�I�[��|�՞�z��֒�k���T����-X��c�m�f�k��x0o�S���7�:��6���l��T��n���*���a�/;��	����-���cp%lJ:�?^|��L�8��ms�|�xǄ���8����$��:��5�6��e������XlO�o3����bz�&�#TLLQZ��؎ɩc�qx��>6?��up�I���t��De������李��zB���?v�n�c��d��"F���S�ÙtU]C��Z$�GlA(:YS�$�v�-��;Э)ԅz[z�:��ԗ)#��(��Sa��ѳ�e ���t�{��\�1� *�҆SR��7Rk��N���pR�N���k�H�ά����6���	&�@0������.����I)�Em�}�#Sr��芗�\	�jh0���1 �+�~G�.�#��ͽT��;���W^���s�눼�c���S�g�Оm��������%��*s6��������#��@eېvl�A�h�;Z��x*�)����@ju����{� �7�{�LI��#�%٫�xAZ[��W�|钌Y��~3�-c�>�_�U����*	]%y�F��Љ���\~�a����ɩ#9�sK���/��u*J"�^�;MQ��rv �ԕo����8"��o�U}*]�PS�� f��G�*�'���0����8��b�l)|ETsiDaJs+H��+��Q�ek��Ԇ�.�~�n�(N�sp1�Η���+��R�D�J����qP�e� ��e?��X0\���%�H�?�S�u�k۔7tkk����o_��O�l����#E]���C�6G�w�/b�������!����G�����٪��W���������w�!T����jzܡZ]99U��Oʢ,��������@����0�6���Di�D� ����+��'	8!����wg���i���}���o]��2p������FiÛոU�O���]�j��%9�������*"�{�ݳ!�WF��Ox�����Yz[G�Z�A�g|�"+\!�|�VA�g�}؍ǹ����\�.�M��Z��M%���>��~��7o��i�)�o2��(��+�^�b%9��{le��"��>�|��<:�����- D�_`g��[����Xj���]vMr�nq(����$5�.0ڛ����D��hrǽ�.�����_�7h�=Q���wilJ`u�8M�z�4��z=���A�{׭G���L�U�}��KZ�S��rX[�&� *��N!Q����&�^�,$��lW.7Ƽ��Uƞ_Ò��Ў�6)/(�}�#�K}����/�to��D
D����'!�@m�<���f�]9z��8x1�]C^�u�^Ep&��k�&<꺢s�\�����9�N�ř�^�i�}�9 ���N[^ ���_���)O�����?�w?�s��Z�+ϯ�&\	�B�i̴02��e@���MB֚m��f\�V&�#m�|�_b���3����m�Ú%^9\|D�c���(l|JS�+�`�����0�����l�@�L`"��]>jHx�)� K6rS��o�wa�w��A�����D��y�����۽
&�	G����m�ݫ��:N6��mM�#][I��j�j�od~�0�QF�)���Ńt��{.힄$�Ŋ0�n�W-bG¾��)wɨ�5\�m�2F�"���N��̘�'2�����i���e=�l�N�ͤx�52ݽ>H ����QY�jG���}�� ���K~�7���ͷ.[��}I?���ؔ���:�n�.�+T*�,��w�ۯ9������%��/+nh�g�ee���4��a'tB�"�/�Z%Z<?�+6�a�����
����vgx�e��� �'dN�K&�Fj�	�E��K�M�J|��O��xq���3AsƬ6��OL���5�
/>u��BT�:���:*��r�o������If�i��s��ځxت�r������Z���vt�!-/�)}�����m.Zbf#ٮ��H+���A�4C�Z.,��'b� Z*W*����E��͞�&��CЕ�Iꓑ�k�~-M���aBN����I�E�)��d���K%2�4tm�B����3\;�/���t(	e�=M���˩!kdX�Mh�Zk������1��j� �U�2:���J�����}��p&4�э ,!fh� HY��Q�z��1�A�ON�ӈ��	�r5AҏUK0���W�+�j�WLr-d�I�?���;�3��؜�o��Ƴ5W�n]������!
���^��$�E�����^U�-6��=�zQ��, O�SG3=h�c����{��{��E ����+�r��;�O�)��C��~�,������Ӽr%s)�<����:]�W^ZV˶��n;����y�u^��/�ftl$ƶϮ�KQv��̣s���>�ѯ��'}��*zQ�2�Nl��+��n���2�����܂�U`-֦���:ʪ�f*z�� ����l���T<�h���Y1.�q�z�󶠷���~��^"#_u��2&7Y�X�6Pł�?4�M�R�@���,'�L�bTb���,�� s~���}˿�]f-63ۥ#7I�.�V_����po�Ǧ,�]��䛠�|�����Ϲ�"��������7�SA:��x�s>7��M)�Ur�����8�����[/�)Ȩ��2op]�e?��\�=�/:���&d��s�`%� /C��0���[)ڛ����1��<B�m�Z�]ה��V:�F�m�������"�~\���;Q���3��|��p��t����e)�j�E�i˳� �8E����8s�_���:�h�ϑy �X�W�چ������
=S�Y>~:�����?�x��@�u��E#T���'���^U����O.�Q5.ț>#:%���4�v�m�]��+�.�[�]K��+7�T�����Jr=��������:�:ý� ����Cן�K�Y��t���X.�G�jr����2�|�o�=p���*6�RG�#/�:Q��!w���%t�ӂ�ڱB���ɥ�Y�CȔ��
�e~I�cw"��8�ꢍkfJQ��Fp��7�fO�>�c)PH󽳠��b/�j���'m�Pp7B��Hj�aML�U����o=��ebEr@x;�cjN�K�'7��j;:���y	^��c�Q�HR=Z�I���g�1��0)p	׍�wT�=�����nAJ�Q�V�n�*55^ǢQ�^X�����N�u^M��g�UŌ���(V��.���דU�^����Nl���v�Ԉsб�Qq���ڽ�^����8���?����.�g�]�l�#���}���Ytc�G�L���~��=Ǥ�6�)B������:�B�9���+�R	QP��&� :}��lHs�!��c�bO�7�PE�$�һ���
扫y���Dӫ��ʄ�`�y(�L�' ��O}���n�����,�hf����g�3$�������a��za��̷EU��i���?�<n��)w����Χ	�q>��ڃc5����^��6���]!-�$\5����i�`�`&��b�9�u��S�|
Þ��V����$A��F��(4	�pTՊ�jn�(�sz��>& �$S�[g2�}HpF��i��n��lx3�ў�O{�2UDJ�V2�$�
t�N<<&�B~�P̼G4U�d	�$a*N�t������u�C��Q�G53�N�P5$��j��s�:�gtp7.�mg`+=-��Z�)e<H��8���Û���M�c^[Ѓ|x�b���42pG�B$���"���\_&u��ܒf�א(���XUT�)�{x5��@	�󥈯���<p�4J�e?�?Ơ�~��&��V��V�>ݑDƯ|��y׬V��M�#�l?��9oi��4���-��
 g�Æ�F�'6�Ϯ�poe[�z_�S�fc��}�s3r�WU��q^W<&;�r�cn�|L<p��~�k�­����/��|�ˮ�$T�5����o��'�a�k������g��<z�ԛ�C3'}���Zi���R4���F����7�g�Ʋ�l���'B8GK?m@V��4���EYh�����Q�V�fl��m�qV���'Ӛ:����OP.K?L�/��W�����J�Q��_c���8p����p� ٬�ߦAO�P�jAv���j�PuO�o��_�D �<�\e}����C��Ɉhq֍�v�Cg*���TG��x��rV�/��Ԯ�Ae	/>�,b��כ�hV,��,Ί�(�dlE�}�ʥ�/��<�0`ep�������	s�_���{���j) �ȠgkT�= ��ĺ�%j�X��w�u�&��^א��;���s���1�Z����Ѣ�\'Ӷן͝�H���2RIO��*�
��̈�˶�5̵�C�֣$8������9��/�Z9!wZR�9 q��+XM�-���sl� ܢ������=�¢9o��ni��g���Zp~yti�p���J %��o�1���ٮ$�Fc�i�g/�8�`�p�z��K�uUX���xC���
�@
����T��CW㶧�1�,���,/a^v�;B�1�l�$�u�R���%/\.=��aw"�JN%��Qn6�~چ�C�1gIU��.$�+y!0�K��NԐG^��`�v�s�K������Z��YSS "2��Aʹ@��C��>�%�:Wٹ�mlI��.�Τ����bG���M�ܖm��[�����e/�s��a�Ӓ����Q��+�nf�KH�K��ѵ�L�u��Y��}l	gXk-��%��D��
n���́�.�y��D��eZ�xJ�����Є,g��!�da��s�Y�o����XDy(@�y�H�8"���f��!��w�Y�Yc8��7W^E� ��?�'H�ǖ	����0��O?�'�x�"���D�M��_JT1\J���#�ޣC>���`�&?�
'�^��CO��\Z���N�Es��Q��&��yp����Uu�)E~�Hp��߰l������B!�A�/%�饥��͇����I�\�~$� �� `�������a��3��x�5�������U�Ѭ��!��6�D�hW�V%0Yz'{X�A�rF��D���V��Ն���uh���4��C��Sg�	3����&Я>-���T��tlS�A���WQӈ���!-V$F�E���&}�/�c���_�Sp�o�X����D����waH��	�����2S�v��3��&�d �e�s{�:y����
;}����"~1V��<�����Q��{�\S��Y��;�]KVQz�v@�-k@M5�5{ �E�V��:�.���m'[Ic4PתC���D�A�R�ᚄ 'b�^t���-d��W'���^�+V�
�R��*^_v&7��-���:{U[n�5T�E0�8�+�g?RX-{�B �lĽ��r�1����D��^�&�]zk�!�U|��C��>�7k�����C�����Y�h��S]���>&��o�$u*�H�~�p��~��.?�k�.��uN`3x���.*��l� �ːWe�R��c��H3�k��	@��1U�!VE�S>�8}_�G��?�t?W�\\�'��I����R6�O�G���:Go�0G���z�>J2�}�|\~~������z5�ŇAo��$���F�5U$-�e�~���-NF�ae��@ۊ!s]�H�D-X�#P �Ic�Ɵ�g`��L�7X�m�<~�镜Ns��pS��׽5{�|��6�pP� ���+��+2W߾�æ��A�%��q��hٝ��!�-4|�v�5�����j��\%em ������cԪ��7�g/��O.�	�"��D��+�O�*ݿl�t�"�v>~cҁ��d��O�)�d8�Puji����?�V}�ۗ<ȴtI6� !P��bl�+�I>�·�䡆��,S��4��޳߱hӻ�rR=G�v�\z�d\��:���#H�������8Y+��}k�� �Ӎ��9ÒZl�t��B��� {-
żF��^�`�Sb�}_�l��.{x�|�g������3F�Ii��z
���I1A!�~�iO�Z6q-��+�/޼�X�-�w��K�R�yp�sh�Ut����|IM���֕�s ��Z=�O�}�D�$�愠g_�ߚ4�I��Y=�m�\̦ƃv$�j��w;&KgX�Y�5�I�� ��M<�W��)�o����+�=�U�qO�	�:s�=_��������&�;}�g��O�Z�GMhe��}�F_��5�dU�Jt���M�`�`Y���"t���B��@��ꑛ�,��,
"v����TH�c�-WE�A�Će���p��^���ǳM%�)ʹ����Q�P���iM��c
Crh�.������֫3�!k�nY �z�&d��nI:���we��$X)B]�����?�"T�bA�����歘��+�Ck��Y��SY�Zݴ�����||��کK��#$�8�s�Y�������U�����"��M�vn)n~�)v�j��3�6&;]T�Q��)b���#%JA3����s�M[&�ټّ��%�C� ��_7����k�.�5Т�)Z���,S��1اw�͖����[�wmd�t6mcgt`���R��U##wpm�)�T^%r��b9t�H���bd�N�I[j��6����T}��w��>�C�Oɥ ��?m[�/ڵ���G�T/�RQujơ�P����儰�"�|�
_���A��A���i1N,*�=4������]���� ofV1{��l�"��q�dK���W��[�$�iL�9�oћ���9�N�9=��������j�{�$�!���ƴ�<�2a���
yÎ��g�l����Ҳ�9"�.P��,��7{+��d.NU������7"ͦ��^"�a�&�-���7�*�\@��imx*��Fx��!��I�	�(Y۳dY��o���!=.4&1�lq�`H�m���qPv�U��v�h#�:���_ڲ�P1>�{ĺ�A������G���ӟ4�t���&p�֕h
��T�A��ln~�sp��\(a���N��ǬƂxp =����U��2G�^���Y��$-���^�I?4�̤c/�BE�̓��o�rV_p��*#
�t$�\�Y�S�nuuzc���y_���8(`��P�8�p]�CrK@N���{/8ޯ�\���=�������o�pB��A�p�wc��+(�x�~;���[�����&�����dRܽU�I���g���h�p��qB�*�k�:iqJN��42�m`����E͹A���f�~N�A�M/x��U�:�]}-������D���H{-� �uH��x�V����͟�,�C88�˝EZU�WXk7���;�BI�`}���eh�rrJ��m�( �k�h��l�y�g�.�0E#�0lם� 7��T���&��O�V�@��`��<]1�?�Y�,ZjE/y���Ar�^�ٷ˸��.xiDunV�Vp��_��S����?��?u�
�F������-����vv���j;<aJ�%��O`�T��%Kg=5~jT����k�ÿ,�4�O�����2���9�������c�1�#S�@@xt:��%F�e����c��P!�Fד��E隌����TcϸFEG���X qց�%mA�w̩���U��:h��'o����1�+K�'���D��������-����u�Y��7-��	��
nj��%t�{~��\lT�[�ty>q!eF�)`X��DD�"�ȸ�2���}������?������X�8��������!����i1���	~8=*,Oq|`]?
�3�en�g�KЙ��(�\'�^ڬґ��
�k��q��>�`�n��]��d`���P����	��d%�=ʩ��VbE���!�pm,�Fv$] ]:���]�dB������7v����Y��u^Ѱ uո�F���A�7���hh��I��P�쀂_XCV�\`�)��{�^�����Ur�Ǝ"����V+3��	���\��`�
��{i>J����.FT�w��$�
2�wU�t�`2���B�+�o܏f��=#���Y���E�s�S��\$kp0�9kZ!�#����܎�Ѳ���
�U��ˉ�� z�@�}�s�s�<})��5@�����ճ�o��%e�T�����5�
��7d�Њ�E��3*Lg��@5{��7�I�R&�7P�K�hݽ���;Fn^�~�su���Le�P}��ax3��,%��W�S�29`{w���T����lZI��݄vzm�%��#��fb$�({���C.�&ג�
jm�W��	Quv�w{�7���[@6׳f�3n80�,�-���U7�&�J�6]H�/�����ޗU���������ɲ�E!�6�J��P6��+��-h��XљnT l���-E|���F�~i�d�;i4L.*����2忌��R�`���t�D�8ܬ�E��[�'�Z��;��v0?���P�Jؘ�\�fq�Ǚ�(=��^gFu��^��\y!k#tc���G�����(�)���Z99�?���K�N6�&��iС/XהQ[��͵�C�=8���O"����q�W��	'K�b(�oa�o�kS�8����b�~^c�q?��eM�8m���[�����5�sP�!�E^Q? K(�L��8h�9&���M���4�L1��u�\��[P2L��Ty���2�@������sR�ll3��;�<���<� |@CňQ���J¦�x��|�i"e��7�&�"�ܬ	�v E�x�(���/ڂzbP�
c�������=�o��Y��Gd�
�N�5�K�����\�p���y�:q]Bj78����/�1$��Dok���Aeן7"��<����W*�){t���s���T/ZHI�ˎ����,�S�͵���K�$�~�:�A�,�%	�C��|�r�!�ٹ1!�Ű��c�4N��j�}�(�[��k:W�[l	�
6��Աa�C�t����=�� 0�)%2�>��X r�E��a�W��Cr��t��-bG��R��Y*�Ӵ��όͬ�.��~��J�[;�����:������C���������<ܩ-���zw��� �Ni��.R�N�d�g�H�k��r>E,��0�YV����}a��r�������
lz���>Ɨ�x���T�5ؠ������Ir��Lρ`S~U��>&V&��Ȅ���%��scf�"vھ����y�|�b�̫U��� XSv��:P]�|:����,�Yg��L���4:`�����B�C>�Q�A����Cа���A� ��7�����ak�U0m*�`���]�ǠmY{u:�����y;LhZxL��
a�C�;rCq� Z{��i+����M9���N����4Myk9<�V�h�f8i�cj8уBx4�>w��,�?�|����!$�_ү�񛙑J�[K�&��D�
 �+BL��ؼ�N(�2�X�p��;
vDKȪ#��u��g(���_���)	��|��iu�wwdZ�B�/@D�J�J��������]�t�d��,2��^�D
�����8�ޭ�K*FB�S� >����1�u"��*���Ѹ���|컳ᴮj\]ù�_ ��vm����@��1b��|� ٬Y�J^㽥K��B���ш$W�������u��n�>·��K������� �!3�<�9��_�,]�Z3�!�M>(����,W�i<�xX���v�yE���|�~��M�~ }�$>2�[��l��}^���J䶞h{*|'\��ǃ4���+�AK�n���Ǥ�����4u�=B��9Ͼ��~k�r1�� 3mu�"��������kܐ��TC^�ט� �e_5GN�.�Ï.G�f��Gvt1�k�p9?�X��x��e��j��dw4�(�O�!�ϻ�P������t�T� [5s~��
+� J��Ug�c=!��:���l7���/ =c�!��G:?<���D���yfE%�'!�Ji����I�2�Ў�Y����V=.s?���3
�!���t����	_�W��h�^٠��@����H��e���l9#"[mH��`%7E�Z�O��}I8�z�x��0xH�Պ1=�M4�ˁG��i���X� 3P\}ߘ��qkt��r3s�=ݞx��@ȼ��S$�tn�̕]��l8�ԝ�p
uU�3"U�#E�F+��/�D/Zrj�E�M4%����Z{n� #ezH�~�Y1�M�8[y��!��4�]a^��ؓ�5��`���F�Iҥm!���Y4�>br%E���I��e�ڌ��N�@<�\����������&w���n�c1���i������$��:��J�c`���Z̋@{8����x��Wi�9��n��ʝiѫ_���n��`2ΧHW~��+zV��M/�M�Щ�O�'J�	���p�d�S���~�]�_�=��2|������N��S���q_j������\������b���;a����P���8�x[]�2�TA�N�7��gɴiZy��y�X^��_���R��D��-Υ#��n����0ۖJ³���WV����˂�O����X����~���z��Gkl���w	/A��}��&��hFaL�o�U
М'�/�_/�;K�Ê��e]藈텧�g���a�P�eF��p�^���:�#3��%�(V܅�ք�׳�7��γ���(@�3��e�y�5��p$9��r�V��o�Ze/�8a��9ǔѿp�j�^ �Ժ�༖G�<X�YK0�`�Z�`���+�����2�������_���pd��=�����cz��;Q Έ@e8T�L��R��x�	迮P���Cn� Z�����~,�%΀�z=ʰ��G�����1*��������Ӄ�꯸9�!���'a�ԏq;��Z�[��8R�(��4��k�ST�9��]�NuX�1�u�HS,���K��H��(��GeW��Ms���}���+��@��+�I&�C�e�2���$�����c.w�aG�A�*�jj�Ϗ?q�j�a~D���'�n7��'���+�L�heB����Hs>�͒ʟ�	i�m:�+�a�o�F��H�:�I~M3��I���Ջ�<+0�N|����2���̴⭙�Z��u*�h�B�J�I﫩B ������f>���Tn�0�t���S�����{�f��g�^�%./z��Д�_�n;�����*p�%|�4�}nteL}�;*������-�t��.��!K�]�'tE%-�������n�~I�j��eZ!�5c�K�H�8y�O������i N��
����@�OV��%i���Ң���X�!W��t�}U�E�F�B�$��C���m�^=�P���	���%��UD�J����$���D$�9�K��*�G��C�ϲ�����ȴb��/1�|��3,��zv�嫛;Q�@�f�B�S�GC�.�	���jҏ��f���{2�%�M������mE���+���!α ��FZ���bµu��(U���o>>�a\t�F����/Po�u��jeR)�gʷ�`>s��Fl<�*Pǁj����1�	�f��/u�͏-���l���4���v�[U���� �,9SW��Jdh�ف��NsI<����$W��#Vp�QBMHu��k�<�%���\�>�#a/�8�s�f������(�R�_R��zJ˴p��z�+Ա��f�47k�Sd�<�˄R*SUQ��ᑷ!!N�����0ZYԇ�U>�!xK��@Q�ZRҗw�B�G,���gD�����z�R��C+'�ŅK���3=k�l%b=9ٰ�5c�J'툨e?y���_2�R������~
D��8�.�OPELx>4xB�A��>Tz;�����aL�h5U���
�bJM��n�Py�y�Nہp(�c�J�@7?~\�F��q�A��i��G|��Fv�K�#N��?Q;�E܋r}���S��Smi��7.JW��m���O:
���2d����҉���[�������V�̴��e9�Y60,�wn`���b��	��m6���(#�.0��q�%�	Z:f<�E��������L����F�qt�5C�2�+  Ӑ�)'P6^W��M��N����6U���N�֤O�"�T�?��~��,HA�����mi��U���4玞��W��6�������(*�<vq]T��B��<�v�w��je�cXk-Ί������0��pj�=�f�����ݷ��o���a��2s�xh���2!�!�c֕�m'��kwE�a����i����(I����SV ���.�S0����B����Ď��p�9tG�m!�X�-��b�<z�����8Р�e��Ƒ�t-�j��z�>�ma��q]��~�u��G�{�b�3$�t�� E��3n��?�4�|�ش�zKU�T֬�Ǒ�DS�Z���`*?&Ad ���K�oG5Zx� �'Rj�H˧Uw�}�0�"��1�Rt���ۡb�Z����{�3>9��r+�z���aWq
YU(�1	�%�������
/\j\���nG?N�P��RS�!"W{[�dd�"U"YmTEꁋ�@3\+k�Zuȸ��4KG̨S�H+��s�����Pc���	5$&ㇴ��j����O���Ȳ	CvQ+� ��;���!m���2<�KT3�p����S*-l�����9�Q��~���qҳx@5hV�E�����_J<��p�<�*�b~���!�y��YMy�+_�m��_��H������`���\���S��2?H��y�`�#���Y��f��i�M�/`]��|�d��5��M����eB�n�:'�c�M��S�cO ��jEN|sivt����O���S��,>4����;�-?~�SH �Hѣׄ5�3a�_��!��[��d� ���|xR�j�Y�.�� ]<v7}�o��M'J����4�~ 5S�� �h��_����AO�F����^����1�Ʊp� _ҍ�{~Վ���=�/�;x��>\a�֭ט?ֆ��E�������q��;G~ݿ�/���e�j�Hx )zP�vZr�U�����X���
4	��}��,J�E��$����<��wE��կ��^E���p��w��(�[��ꯦ�@5���B`_Z_� #w�F�C�V����t@��S��4�5�n%/��l<{�mk�f#0U���.8��!	!l���ҩ�w,�R�$�)K^@��s$Y�LGH�_�����|��_���u�a���z�==�+I��!��L�yG�g�O�oN���	�P�H������@Awi���e/]��WT�t���E�k��"=a&J��h	���M�Pe�	�U��V�1��gE
1f�Č#�zϱ�`ձ"0�8�/L���q��:�iL*��v���P��G����������%y@���|.�t�*g�V�3�:Ѯ�\thn�I��k5����u�Q��)j�v���!ICݞ:F2+k�u�GR��@��V=/��ʘ�70��7O�e����@$!1�!�r�Px4�4����\��>zS���T��.�g�=l����˳�׾xe󓟐
����48��\P��NF��9����zCbQ���a��e@�~1��(&�s��t.L�ͥyo2��ISܜ)%��w��}��y�$�c8�>�/y��)e�j�O�C�P�i���qvN�AB�y��w�p�QCW�Pֱ��l�y�E�%D�(�ǑY�+��s��>�i�����;�O#VzVOis������H�O�i�����LR��i�R�$f��2�O��0S%��2be�%3򝞩lF�ی�p-�U�p�/���^�OE͟�0?���AA�%B8,�߽��*A`v�E���@)��)��.OY��i��K��X���OE�j�.�������a%^��-��#�i����j�7u/'Dmjs�=�pմ5�I�eփR�B9l���D]� QB|`�y�l�}q^���h�)��_���w��/���5��Q�~������$�SKֳ��t=ʟ,+t�"hu��@�h�:��2;�ߋa�
���܀OΪ��£�	�ȩ�\���F{E�'�r�����G��:-֮]�dz̓�Y�V!�_Ef&=ޝ:���x�"��O��P�Ð�x¡B����`J>Nw�B�p\E���Ц�;���C�Ϡ��sT��B�,���͒��Q��/~�U#���&glz���\5C���e��r*)�,6��\���L�e&ͩ��\
\+-��e�=:�Б�z�	��v��j{�R�a��BF���-pOcA
�A`����,L��ev|w��d��Q8��#��EF]���aHwޕ+�c���v��s���BF�P�F�2���ڨ��$�94��t�S�n�(�cKT�]��Ka������J�s9��FV����PX��=�ƚ {U�GG�x�UC�DNI'*�~��b�������ί���Mv!Fٲ*Q,�}�$��ہQ�g���irw�J�F��V�"N)	�HR�9GT0�@�Q+��)x 3]��Z;����}�x�}lw���L��՛�G1�2������N�ͣ[_��gK��h7V�=���V̄*����3���3
 2�`����Z D���CR��su�5�����#�.��+=0 ��``�P��e:	��>X���J*�	���܆�s����8� Aa���a�t��R��7�I%��m���zH��O�EZ��������y�a�8Z>���v�h
�l�0Dk�����0￥r��+o�o����F����Qf��	��t����NWI�%�l_�Z���.z�2o�lL^����=��A�J?���v�[(|��,�t�8�(~����>H:�n��B:����㵀~Mf4��R��&�-og����8)ڌk^S6C(Rʠ�{��6���E�J����#��.Ɖ;���
Z����Wd��yژ v���Xߏ���O�^�<mF�J����
����5\�����L��-�",Sc�?0�Լwdi�}h����6{��Õޥȋ�
���ߜ`g*�bΣ�d�k.��A�9b� -��\�^;�/t�R^f�\_�����
_��!t���3�q�	C�����N��H�4��վ��m�FZ��M�JL�A�l�4��4�1�IpN�ˏ)�sY�3�A�"[�q.@�։�<��W(#tN� �ݻ)��~�J��5s�?>ByT9![�n�)w[��,��ݙ���zp����_�5�� p��8��-z��r��jB��N��NpN�R[�K���x��`&�+�Wv��ֳ&���)���չ�Ŧ��;�41�Oc�hl~Z�����X��_
�4\��}��U�FV&�c�q�
2���,��n�4�����y�����5����x�(�#P�A��6H����H�X>�9�!o��|$H��ۙi(8\�ɍ?��G%й*�?{p
�$&���(`<Ѐǖ��Ě�'8u�꯯�-�ѣ,<�;���ކ���bd4�K�-.�I��*�a�Ǒ����a�^��Q̐H��ch��:�8���('�_������$j^��X�(gJ�����r�V[�c��dL�K��c�	�`�j�g!����s�bQ����2�W��S�,��i�l�i���:0��Z�'�
0���A���Ƹ�)\�C�,�E� 6��d���˯0y;ͦ���?Ӭ0^�XpQg9r�l �zТ�(h.��Z��UA��[4&���§1��% �5����*�eؽ݊-�^ѭ��{#�9�䔮TW��_��GU\�^{�F���~�4��c���������xN��A�v���3����VW�<%�P��3�h�XW���ae���36��vt(y���YOUPAr���W��֛u�6ql(��D3IAo"��W±��G�^1kE��x�;�q��_.�b�<?��aX!՚;/����Z���^=m�'>At$)5��]Բ�?�#m�����栧�X���/+,_%"�c\>��&��X�! 1 ��cE3C"��'E^,�v��5��f�x������q�4��,_uy�T�&Oz�@��Jf��9�%�����FKD}���"?��9�����m���y��H�I����pM��dmc�E�Z@`r^�U���mM��Om�0F�{c��y�\��K8�`�b`	i�5gPQ��������O߭�7���������Dî���� j�Ձ3��Q�|B�ɉ\�����.A�A>���d�`�5���A�Hu�G6�CԸ��)h�3}�r�����S�nֿA���I�浪�ܠ>uI&n����M��t��7���_��PQR�:�����9���`�#8��%��A���;�N�0�s�ӆ�V<����5|����.6�v�j�	���:�d̫� ��K�l1@�Ah
�4�"�.�'}�ŅyhPAd9�y5SMu �c� �?d� �8���@7�ܔ�H�`�[Z����`��@9����R�3$�T��K#oA�B[��^n��YY��>��y3
ӥ�����oo;.:����x1!t�*¼CaJ�߭~}�mû�J���KyB4"�:V���xR���5]������jOj@PԜU[,�\n^�E�_��_������6Q�D�R�p�!��x]��9������EbCP���zj���(�&�_-�k���	&��JA�=9f 
sh�gLm�+�W[;��J���&����B��M�J$vj����r��b�{�K�ĐZ�'ũ���s:�IRAZ񈻲jz������|�n����0���'c�_$욄3�>�qs�$�0�3�Mb)�BdJ��w��>�'d�k':Z<'� �JGƖ�lD��9[r�i�IX�A����,�f-��t�ի�J} &E�H��K�.��C���%�����d����d�J���$Ah �D�!6�
��UDy��yB�g+R�'����{��j�#��#:��M1J�G��8+��-�w@�a�أ�Y�)R��غ �	�g"V��W�A������>��,3Ǉ&V;f1o�5�(��g�[N�Ǩ-5b&e���8�EA�G�y�jD��_�ѕnq�(�O�� E�o��^a�A�7ʜ�F�%� �v��˝�E׭aԀ��;�r$S1�-O`��y3��i~Kn�j����6��B�ua-a��F�in-h�QO�[���VS�!$�wy��p}l�oS������7Z���tJ��*!5����ǩ�?Np�>��I�,I�+�q���:�#�"��_�{�r�&�J{��+�˗��3c�A�w�T�s�,X^5���&�2�N�$0zI`�&�VG0�F��*��c�HA�����,���4I���s�EL"�������̍�U�;�N�Uu��8
6͏���,�t�aJAO.Ώ�ɩ��%�l��!�9dlj�H�����ق��f�b��B#uW�����D�M�:�>� �Yx��J̱�^$�/ȋ�uV���](���(��=@��X(��B�m?6�ݻ���7*a�o�L��gX���W$俋Ye<y-�n�|y�&��*U����E�)�+�;x��YG�\�����p)�v��F�v
7�!Y��jd�)~��̱G�M%�n� <~(hcKk�_+$v���I�]��\�G���I�h�����>Q��Z����K�4*F��}]^��S���e�K�n�,����=]Y�ѩ��X)�,��C����M̿	�5��7@�3>���b��Ee!䔅�YK=�-	t�R
�ZxOzlk�l�J�*Kk�keʙz���c:�#�-�艫|��c� Ÿ��J�i)祶���S�Y�Ϥ
NHY�Vuv��V�O�E�-iV�W���M�qU�nf��k�b��8���?�H�y�
]_������s�\��g��
P�TÑ����I�Y�fj.�������!���EjvE�h��j4�g�12��i���r�\��g(yBo򽍼���WJ+z(3D�F:g\�f��7�lҥxX��~.�_����t��Re�=�{?�YH���`M�޻��)�