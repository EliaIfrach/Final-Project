��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��-�ro��i�����/L-�U��lOjj�l]I߫�p3^������_"�'j�ʬn�*W�� �a��;��}���������)t�X�|�r|�~U���;��k��2��%�`�	�c͜��d����/�OB��*$�K�[�>�)v���������~$�sF�]����ZP�6͝*����ĩ�';ɒr����YU�|��#��Yq���65��~�Mduث6z\j���4���E_w3�Cن̷����o�I��Ƃ�G���~T�VO|�θ.YW�9�����I�0�J����r�=fw 	`2K�$]�NF^-F{Ux��L.2OP&~����k2���S�BY�F���iG�H�E��+�%h�<����I�[��G/*/�F��➳��nZ�W����Y�o~r��_�$��\����f�M8D�o�OO���"��D�_U�@��MC�`��.4W��ف�O(��
��,-�h��jn<;���#��'>�鑩�!i����8�1	ZB4J�yY����p>G�����ٯ�`����?C��?��=Y%!��b�IWx+����Q�XjD�I��5��� \�u�u�@n�X�gs"ݚ�i\�X�8�xt���'� �� ��\U,��P>�Q}�������g�]�JJM,��𺪆l�
��z�G�+�QeE"�<���?�PS��"V������FSh�Q��p!�o���M|ln�P2଑��\v����7��e5h����p�C�M"�-�v��4͵ȁF[�=0�$^��ܜ���y��Q$u$���6d�
��"Ｚ#�/��/���34�}��$3#|���2���"�f�4!��Bˢ�mn@��Q!5���SU=��h��qJMr8�q�<l)�Y��Ѐ��������eg�fMV��I-iҷ~$���^e%�����^?⬄�٫%����@(GI��}],#&�]jY��?�����폿�����g�Z�+	]�Ei>�X��0�ݙ�Y����s������]'��Hq�M��B#��o�9����g�fuJ�b�Z�$�Fe�h��<�%���Ȥ��E��x��ӓ�^�)���H�^���`k�2����IZy��%�AO��b�}jS�tX�r�M�a��6�/e�/�{��������4�l��A�9p�P�!l��?4�)r��L]ʨ��?������ϚYCzS���8h�,�5QeۛF���!� �XP�Bɞ���m��&�z ���т�ܸ��2Hk3���DEM�I�P���Rtn�9W~u�{b9�\�E�Z��@ڇ��������^p����b��Y�N�GǗ�ֻ9�嗛rWQV��},#� `����S.��dL��u祥!8�����K��7Z����>uf,��A���W�y�_N8`�|�=�CZ����QHu��{u���6v�͍���w��"�~�$<ݬ�ߓ���@�C��V�$�E�ү#ڶ��W�h��6݄٫�i@���u0�E�<]��]������D��7��e�C�s���X�.&�@����׉l�X-���� �{��*�S��-~-�5�H���0Ou?�h�T�p��Bh���:��v�X�]p� ����e���� ���m�k�'%~�a��M��7�hʅ��U�Y1��Oe�`W��5��j�����QS��lP��xG��[O�}w��#=L�M�90S0�r�
��LX����=ŒCZ�+H��-C��8�0�����z�m��Tlǋ9Y��l��߻�}�7tǚG�vo9PO�$I�@�N���ONj����
�x?�ۙ#�##�n�y
:��^8'�X�0L#�Ş�L���A��S��K4��b��{�\ k�H�M�MʘG�1���+��#o�[Jo���A����7Pr�Pg��N�
c����E tmU�!c2>Ԉ�ݵ���N�6�N��~�
=�ٌ��TרT�w��<��ƅމ��6�&\�P�@�"�����e�t�� �X$8��T|���i0��4��;�%یvH�����'Pt8��Ns����<Yvq'b���Ǥ���@;�YAqw�@��/]�wn/
�M����X�*�N��(���ۼ�HHp��\2�=.���jmQFs"}du�-!�ރt�`^���H���l��u�D��bH���;!sl�_OW��kO�F�w�p���8Y�� 0[&������q�O-n�QC�GQB�~-��M狅@�Q�z�.�0,ѭh���49�ҖO�N2�=�
�o��q�e!<D��SJ/<��O�qF-�{��Ś��§�>p!��M��K��� �qFt4\�����0u�j�H�$O�{��9���CҖ��X~��d<��-k&�B��V�r��ء8#�?�R���c�{g� ����'����m�,���H��7��n6̑�P�����7ӇN�g,���p/���������a�k���	_�h�|�Sq��w�}�8�Ik�gk;5	O�x�h׽�+��������0��a4{!�M[&F�{�Ke_d��jN���|:������<'���j�^y�*��h}���+^ܔt�񓿩�F/9�ea��&�����9mh�u�:L�9�ʎ1��d�ҹa¤iw����9F{�R�qlT�)$m� #�^���� D��p����eKڌx���Wv��7�<���Z 4��d!{]'+nJ�����7�c�V�%��s�@�Hp�ƊO!�3�W.�-؊�<����QK�XFs�'��x
i��7���iyx�	D}�ɭ.�j�B,�]^�a����p�G�a��g䬗�3-R;%����ֈ���@�v(<#����3a��\ �'y����廛�5JbSl��E4�&W����8#u�f>q��q�MhZ�g/]rm��2�?8b��|��hEq�Wc����ʓO���]Ƞ�٫p)M��[;��nO���eaub	���8�[�%�m�?��!|���>L�~�=���Efϰ���K1Ӊ�ך�	��	���b��B��O
$��۽��0۰Z���Tx�P�O���ġP��V�Ӹ�9g���ϩ��#]�1�TבS��������)+js��-�[�}&��V�!wZ�#��b��5�|�u=��;n�;�ǥ��Y�Q�7e�3��ٯ����uy�K߰�f�s2	*��kO�_�U_��ե�2�Z+���H�&3�'���x�0f��Mr�vb�ZN���h�kk����FS�0���	wK!�p�F�EC�(!@�O;l���Q�-�g��^�U�}�Ȭ�p~A�D�/����ɥ]�S�7f��W5��[}