��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S�OO�$����d}�嘩q7� <���L���������w�Q��|�7*)⠠���Hf�(�Vӗ�����؏���M�(˔�Ywm���"jN^r�Wf�k[���_�)�q�[ţ��!�&� t�U�ܢ����G>)��vL?{�k����Ғ4�1���%�� 9�F,2��4�"c�<�:ϧ���Q�*�p�M�^DV���<��(^����RU������xS���}����m�����,���kCc��iE<��	�*�t�c6�2���{,��h [��O�5oU�!8�i�S��R�h/���"�$�sx*Ot�k\��!�vL��"���+N6�>e��	�=���)j���&�|`'��2�����ǎf�� ���[����%l�Xﺝ�:R�V�m�ɧ��;���w��ռ�Ï�;q�F�	��\t;	��6 �V>˛ߟ�oGp5��-���:�2w�|ʤs���D����tL�4#�o߷�:�S�|�Ȑz�C-(�=��"�4� ����F�M%�兓t��zñ7���[����q��(/����M��֨&/����\���\�&�d	�� s�% �z��щEg�pH�eQ��#0�mG#xV���g��I'gIV���T��B`$�\A�-3Y�=���äJ޻WA����nA�pC��+2�"��l�����7��_���������0^���uO=�̖���4����`�Y�v��W�g@�kP%����\t�
��n#�c"��@���o���?�z-ɐڐ� �ȇ2�O�U|���J�;	������$b�,�E����E�%_z���{�GB�g�����֠3r�؄q��lX9�X�!�R��h��Q�	�W���כ���w�����8�]�8�ׁ"&u�� p�.�Ϻ�-.���j1��vo��r��	\��`ܣ#�0��'��tq�Yj�C�I] I�9*m
�2�\LD���Cb���T�ä�y�֎{x��b'���:����U����o���r���Y�$8�-���\|P��n�HH}t��2=N�˧¼�^��J��2.�ǽʔG�_� c���t��8)�1J�Ni���<��6P$�T8P@����ß�����g2���T��z�L�% |7�:���?n�Sb	�d.�~�W��^1"f!��]A�p���?|�m�����+5�?��ɔ��	Rdѫ���r��TC�:M:��{2%Q�����uv�/�wk-'Z-���IU�Q%O��Y�����BE��a?�'a.�� �mz.��6 �yTi�~:���%�N�Nr���eh��sd�^�V���a n ���ڮ(OZ��\茖�#�� �(���S �e@���?9ָ�w�O��fN[8=M�S�P̻$5�r+7~
|�m2�����E��|&��js}DV��Ô��ɿ��M�3mлd�LU�+��L��;@�0pi�5��<KX���g����HO:�[�}.��
�	
d���qᅺ���2�Va�F�DS���2N>)�(A�J+{3�FE�!����h��)%�����w�nX�+g���$8�=C�F���������G /ZnNS��a�A��|�6�)�r,�b�����ս�4c�Nh�����Lq����Yecm�['mip<f�C�tν��G����p���z����:�Z/Ծ�s��"����V�������F��Չ]���J���~ދ �Ȯ�0m�#�H7sP~�4��p^
)!q[��&�ްy��2���u�9աQg�`��8+�	%���q��-0w7�4J/�ͱo� �j��On��F�FY"
��:g
�AY[[��2�0j�ʌU-3T��������~����"��2*�{�܎D�W������%�6eFFHB��و��$S���g��ʊ��#�|��T+y/Um����h�aǁc��+c"��&l���@�$!�2A4��Ř�Z�������{�[�KU5μf �jm������� �� 8�l��cS�`*ϏZ���&�O�΀ ���Ri�N�",��G>:oïc���0�^zsɁ��+)� �em�wC49��c�y0�)��d6[ܜ)�xu�{PMk�&tfl�64b�D^�EEw��{�:���G����M���	�e���H��s fo�*�*��Y�rgtI�����>_ĻF1R��U렊:���6x���30�mֶu�C.t�	��[��y����Pd�'#�J�5��X.��>��_�XvF�����h�zE����5�%�
+�A��ʜ���b`7�q+��?��7�1��uJ�uq��3�����Z?��7w���C�B�s˿W�����	�29b�QQuw�aN[c�~E�~���-���x0P�鋡���
S�a�h�}N ��3Ԯ�ۻ��o�	J/��kt�?�~)#�ȋ��W�WQ�vM=<n���w���$ ]<*�ㆌ��52���"��/��<��@�SQ�g7fuC�e�44�Z�-G��Qr5�1}i���d˳d�����<>��]�q�B�>��m����=���g�u��J��x����I�K8����[�/���k懭�@c'i��޵$�������,I�0��}�+�7J����ֲNގM'W��S��y�ą��D�3#[ʭ��t��4�g��d���hM:z�?�_�-Ϲ�3�ӵ8�@�# (�N[
�ٝ"Ѓ�2�э��z&?=>��l�p���9�R���7 ���{����#��fI�]�S�}W�MG����=Z�dq��.΁cǂȧ����G�۫�.�������s���B���3M�DX�m[:[�~a3Ux�1��S�/Q�H���0aA������?·�B?��A�T��]WBM�W�@]X{h�������m$;̲y�߬�*��/Gm3��.M��
����ֻ��k@2�%�n,����~�VP?�^OT�/�bq�����x�<��:�t�]�g5����!�YP@�>������Lj�,V�<� ���ВiEU����߆��C�b�i9���YyҠ�o��c�����}ĊK3�Mxm�k�DU?n��i�S�
�-/ϒʃix6M��p��͕��>����j�#D��daޗqi@�98AД��>�5e����ی�	�XӮq���uTɃ����e��d�&�H^ۆ�� á�d*񟮵0��$������G���ь�㶪fys���0r	>��
9�n���t�o(���3I�YB+'�ֲ�*��t�2���c���I�7ݽ�������"q#�Ni�p��R��
y��l���Z�*�1���~�������Y�LKG�� �6>cd������ޚ��#����af��� �%�f�0/~�@�!Z��s��M'�%,���y���tJ��qn<mO{���2V�X�+	��-��9���r����U߉jb@R1>{��uvW��&�[(�PWrw'n䐪s|��ӭ�Q8�1Dh.�;�2�F�-��(�,^�/4�&wB��B�	gVy��
�(�Fk�?�NV$7�$��dCA��E�m1��E��P-�N��E�Y;>^��#�_�pa5E�u�|��������������Zh�c�V�Tض�k�s���fr�b�B��:�2�*��{o�۷
'��so֧��M��/���.��E���kfh�$�����&��ٲ]�=��ۜ����?,8t�ݛ��=�������� �qKԢ	�p�,6K�?Y�_���ѝ�'�+�O_9����x	CQ������^��U��w.�d<��z�N���8�5��E<��y�L�H	����Ƈ�q�N�M"p5��H*'"��o�a)f7�!���z�|~�`�י+{�8���,k��T�Ӧ�B��Z�r����e ��<�m��=F2BQ�2��4Rs��f
������\n��J���A��/'�G�ӡ���������p���v�Ԃ��wȨ!^0�S�H�#㿎��y[��fc��4e�KuRsA��K.E�(xzO ����p�=H�1T�^\���<8�����R������m]B�1C?ݎ�K�<�-g�W����Wt5jIf|�����\Y��hX�グ�<��.$��h\&��v�?PQYԎ�$����x..ĭ�_qY+�]���f"�ץ��f����tA��~���yAQ�Dqϝ��BW���k�Mv��/���*�*Ֆ�&4u8nb��8ala@�ʅ=Ѩ�p<B7�;�F�*��))�L$z#�|����l���q�\��3�Fp"��%�4ڥ�lom�dU��He
���?�Y�)y�`�3ݟ�$�]m`������G��{"��$��ț�+eө���H�P��x�����WH���h<�g�aXm'�J��2�|��?	�2 �d�ߨ�����KhD5)n�|���kI�����}��0^Z����ɻU�a�����}�T�*����H֖@�n݌���>L�M��^C	J��>ߦ���8iȋ�����ä�.if{X�K�[��P�_d�wS�қQ���1�k�i��`�)͎�OcK�YqT� j��Q�j�P�u�Z��#�MFQ����`���8Ȝ�@�7�9l�[�l{��,wM�u��:���)��x#�����	)��� ��r�6��1�����by��*=6K��6aW���
�S�X��u�eW�G��g��s"7v~���Ԁ�i�C �?�R6I|�L�����Wx:T`Oz�s�Y-��� 8�Z��Vy-���&<:1��t`���S�/?�j{z��%q��"	2l`Ա�fw!9��J�R�����m+ėm��n��M����JP���'�o�A�m�9�@�d�v�?�컢�Z!x�����P�=��7"��8�n7O:D�����Ȉ46�	H�hZ10��I&b�O�a$��VV�^� �a.?$�_�v%Ԧ��ju���5���������4V]�\���&��%�t��߲��x./1L!��فJo K�T�G���~E�r�+|�EB|l<^.��I�q��:N��x-���\c.\�Ell���{�D�F�p=º�v��a����GN�bM)J�K�u<�w��4��&D���o7�|X/�,���]���.��}#���i����Q���� ��Õ��H�";'�TE9�#�ǯ�Hח�!n�� l6e2dw�@^�-��A�V_C�)gV������"��0̯]c����X�C�Ìp��QQviQѬ�דA����^ C͵� �l���Y[��~N�=��Ýu��(Vp�J�{���8h���-��?�Ί{�����CD�Vo�	
��������7�Tv֫�8�|>]�^Ǯa�s�$���D�k��8�k�o	慭w�u�Z��n���:/
6nw�[q�yk�W������<+���� *�zL\�U��KeD�Q�2������U�]��ŔQ�ph��f��Ժ��g���7+�T#9�c�
bR�,O+n"c�7aKq����)�~)k���I֡AY�P�֗#������}�j�!�"!�Y��C�A~����E"�JN˲�����B +Z�Ҕ�#���E�%�qhF��X�)��RN�k(H8"H;��f*�B�(L�U~v�W^����N�eU�2�Ja�[}0�ŅND���ֆmt<m��>"��$D�D�9|����.j:����f�?�@����`������`�DKܖ����q�~<ه��ӷ���e�QŁ9�6_�I�Ⱥ޲�D���yD�lE��oEE%:?�	�3�Z�
U�|^9*��f���Y�O����V)��&'���L�3�q$�.�K��&G,��P���|�����(+TuuN���6��)^�}�|u4H��S$�n�7��|����;ݟҔ���%�V�쩬��實.�Vu��:?��&�b��~�7#�k�X�1��D�ߤ��?��v]���~w�����ga>)��^A[Bl���[���4S��9V<��D�Z̲����N%�����J��O�
��E�W��6��$=�l��Y���I�b�ag�)�����Ir�S���E�H�A
h���
h�>���L��4�������	�C���ҁ�&��n�̘͗}��{�~���`�����A�J�a�3���R�b��X�ՙ+��=$G�q��Ѹz�"gҚ'�U����,#	+R풞&�ϸ��q'
 �}[�aB����ۃ����5h�,Az���c���A�����@ ,ߗ{���?
p�*#ts�Q���#�5����p����o9����iQ���2��w��ꢋ^b���Q�`�H@c�_�>���J�ȣ��&{^( ���:�=/�՝�r��O��|�C�����<j:��{e�˯w��͹�M���'�ص2� c�����<��DOW���jc"�zl�VX���?�0��y��h���)��xS|Zt���ջ딱���� "�7j>�P�Ҍ��#��#��s改Fv�}!�c�R�+vN�Þ����,�*�L�$�#@��ލ1��>�W�B�i�� �p1��,Ӗ�]L��y�d�'�V�!A|4���t����jd��oT�~N��7@�.�X�a���� ?*��V@"�.M7�,C���b��G��}��.nR'�3�j޴A�����;��tD��&1)��4�O�
�o-�t�	y1�1eeN8ޔ��!x}p��;)C{����.,�
yL	����7E��.m�:�ӽ�:TH�����ͻ:3�d��(q��р��tD<U��`G//1��6PS�μ�L��y�БJH���4誢Xkk_>H~+�S[�)��:�@SPt
>���B�s�&S@j�&BaH���;��w#ɭ����&�� ��(�H�s���ҙ%�n�3L}���9�|^�ub ��2Q/٣��Ϣ<c�f�5�Y�|N�R��}��V��T=6��R2��˓o�j��6��?��8B���LIu--���M��ܰ��.�R�k��}�����D:R��Fc��$��psg"���)_�y�o�fg���1�U�F��c�4�iN�o9� :S�+�" $28��Z!j�V�����c0��K�����݌���f�g�,�<��+\�d,�Vb�IY,6(RQ�D�p���T��Aa������14�FBǏ�zn�z'f�ޭ�"��A�{�5�9�X]����d� �3�x�EҶ�O�0��.��ao�D@��aI��;���rS�3XŌ�

�e|��䜸!�S/��5��\5������`�g�a��hXɘ��E�y��U�g���^���ѱ\�<P��=t[�m_C��e/��܆ߤ��ș��īr��������
q�����9�["{`��R~��ٺ=`��Hا�/\�e��Ju�g�6� h�m�o����IJ�_X�����>{�ѭ�]rL^��t��gjV�ᗢf�@�\0�e6D*'���SG��hB����@3�(�!��r`w��m��| |�1�n<�HWռp����$��D7�=�_i�k��gr��韑�^�/��Z�bݣ�.����V,��I�VI)�r�	�9pWn���X�sG�n����M�E�"��w|P=�>��6y���N7R��w�����S��ϖ'�OB
Kz,�M��rMͱ�rW�%��F���k#1!{`2�Y���;�(�U\����b	���Ko�0_�O��o8���}��܆L@�(R���(
�U85Wa]ݚ����:$�Qc��jF�.G ش�z���N�7w1!��x��}�J'jk�*T�׳p_�S�K�����j�_F��8,s	�@w9i�-�6���{/�A�?J��P��q�;j��������8�{ �e9j�3e¬	6��D�sT?�q=]#��oS�pfV(sp�Z�VBH�/�ˇ������u��`��7T�}���I@�5����rL��N�/�����'`�y�JF�a08ϭ�k�_f]�9��n�iu������A�ݒ�<����\��B��ŋU��vN��������w�越�k�QEӖh��k�+(���D�����V�X�?V�����P�Ja�m	�	�<���P�P͍��#t�mj~{?i��dJP�[�����<XPŎ\�j��X2���02��A��-���'��=����ZD��xP�G�}j�aWel�(_����{�<ySIE�X��JJ}�	��~�TƔ:2� l't{X�ٝx;����W#�a�u�#�W<�T"m-'�m�b#��Yy=�q����d\�=��?a�4����/�K���w,S����j`=��1B���ўTG�E±����7�l�eՁ۱�u_�QTqeOGI�9ٙT��
�{߲O�祎���w$���x��Q��W�w�(X��������~�ۓ�9�&�d�l���E>ٞ~n��"�x��j��Ɉ8er�f	q+�����v�a>��AJEi߿n�Ci���n���<���Pfq�j��g㰮�m� 6�}�\MM�d]@پu���Ru��f<��%p����x� ������i��Kx� ��N_A��Ϫ����>��s��[+MD�քWyz�`����В�$��p�����щ̀�Q��b��;�=�qb��CO���B�Z=�8�$���2!G�v�^-*�[�p_��AI�N�7�9]@꫽߃���b4�� ufZ����K���9���8��KJ��T��&\�e�$Ac[��6j�(^@#'���M���j|��%N6�p"_���+�V�\~�����������7��x(�kM�u�v�#̝+tW���g�l$2�o��.4��O���C���OEK��R�K\) �PG�d��=�(����m	�[hn��a�8�ŏ_��.7���}|a��O:Et�YU�#Z6AZZ	x�9��7��gp��DV(jkTS�u
M�4��tx�����ڇn:t_-YR����&!WgӃ�
�ht��V^��_7����g��Gd|���gX�t �&ޭJg�^�w�=^C��A�RAo}̦ug�!U�J>�h���Z����+�u��d�=w2k0n��6
�;���ۛ ��JE�#]�Ԉ����KZ���x#6�1��V"��ռ1�_�fN���?k�__��[Xh����:�� ҃�Pn�̏�Q��ff%�U�g��N9l�bڮ�*N�a�J棋C�>�j�qW���?�hUK��؞m�r٢*�u���&GDpz]�D����ڵ��A<��XB;3��1o��f�e�zL3��Ы^��.�K������Ur��4l�D���;XV8�!����?�����v/���ұ�<�ý$+�P��������=�����c��F639�b���&"R��w��l34cx�?�SEaAU41`� ��,�مD�#��|�H>���������7bX��K�
2�ʸ�\�N�v��Y.���`��B\6ط p�*iqI��ͨ5-1�\�B@��5��mx;���{��M��Dzqj)��$��N=���_k�6R"�����7��lW�@��]J��o�$������
L��ݛ�h@�ˋ�3Ք,j:�0���T��p�%Č�A�^�ɪW��j���'�i�'�;��E(�]ܐ���WF���r�cS�4��)q-�IR���e�"9=��7���R.���B��&�1�Yֽ���@�GsS��F��in���G�Uƥs~��Iec���<�Y,8�#�:{�,k�vd�����-I�ڮ�d:a��_bn������<�\7N����q�/��8��K����r�,�3�$�
�]�m"~l|��3=[���S}XG��_��ka7M�%�nɂ������V�PD*�cۋ��p���1��XS��t]A�,����ge7�"���Ҁ�!��gM
��vl�4��;v&��mѨ]I��U'��ݤ4ޮX���nI���Z̒�n�L۠�9��u*D�R�S�svrv|s����Y3��ռ�z����x΢�G��̍��q�o���v6�A*�Y<*��~��Z�vm���`�j��(S�g���:�zT��u}�O�v"�ll�|�_�H*&��Z׹�T#��m��/�Wь \������3!oz����2E��ì������%�_"6��&��feBH�I�|�:��d���?"��_N��F�h=���9f�օ>�*�	�@"��)G=0X;<15l���V�����bJ qk�r�$�� "s0Jq ܫ���'����3,�8�8UhK��R贔��z�X�3��������=?RN�c�J����2��"G�{U�Z�I�([�U�H�<�	m��aE<O~k���!c��.���
��8���f̕�Y���5u��.�i��̧Dk�`?��Z�v:p�k�?E4H��J�W[�`���>�#�`��k�:�s�#�kp�{�xjإ����=�[�h�����7��J�KTȫf�Ho�����Ϊ�W����c $�"ޖ��Y��\�qva��u���oΥj����L�d��-
�c�(pD,x�x��$lr�4��X*¡iF]N�	Cy��Anf���5�\���>�{�-���h[���Q�z��E  �%/J���>�: �:�4��>.��9�Ь�_����|�ζ��l�y�\�^�lAsZg��H��f��K	�J��܀Ǉ�����3Xv�e�L52wYE�R=�~�,�o8���S{�K�L��ri2A�� >�ɾ�����L��l�Rc���$�8QG�iA��Ӵʯ�He���HȻHR��nmAj��������Ut�~���p�qR��r�'�m>!�֏z�B��43<N|�����O���+�x�B��RnVmsgiֈhuq�ǜ��e!P����BY$IM0z	� ����(r-A2��g��
J������t��Y���4�Ya����s)��w���Q����c4:���pU���Z�T� �J)�7 �%ǂc���b�'nP��W�@��5.�8�z~����F=M^< ��Z��d�e�6�S�>(�9�o�&�aϨ�eb����Y��f�/w(��&aʰHe�݅5�Ķ^;�uI���'�uz4~�f0W��L|F�]�=^E;�z6��v2睛E������L�=����,�3N�XQ&�M���\�݅#f�>�-�Q�;��k���_]I̟����Z�Ƌ��	AX�i�3s����ǆ��L���b�j4�j� $}�9��$�+��|ήT�c?F�Þ� "�m���?a�i�Y������`��_1[P�M�-}"�����9��>D��5[`�w	㊱JU�yZM3�i�͍���pH��%�;hv����l&�
��R����Z=� 	�Rb�f����9/�_���Ǐ��SQaf��լ�%M���	ߠt̔��X�"��L�*��Jhᖳ������H]��I�C����u�<�K�Ɗ�")%����4>�U#��$Vl�-�f��^mT8�iR·��L_Y=��l�!(���wm7���B��*.�����_�x�qd��p���Sp�dM��,']u����7�vƶF���"��}�f��=y��<"<��1�~�h�m���)e)	~v�H�׏_t|� wC*ʠқ�+�ULx)�;>k�~2P�h�l�3LO�{�2͉A ��9��g ���[��G����i�TK���>p�4���U�T>(���Ф�ݐA��;�@����2ǳo��8\��}�A]����3���R��3Te�rc}�M���
'�'�߹Ss|��9
�B���s\�*2�8��������j��yħ)9��#�>��Xf]�;�	1Ъ&z�D��M�e5�������$�z����y�`ɀLҳ�q�F|�=��Hĵ^�m��\fA��,���[X5��;<5�kP�Wc��9Y;G$���
'�:���� v�pH�|#2��Vvאָ'Vw�0�,贸��