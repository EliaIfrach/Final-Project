��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��dRaXk�l�����>����M�t� "��I�f��Z(|*��h���n�������*)�m��Ha�:?����Y���(�aӞ���!a��,���y�*�FM�] �f�p~�{�
����ז����>�AoW�(��}P$�7䂽�u���}�Z�Wx��b�8-�����J�_]�	@7_����z�Lp�6�bڴ����B~E�Z��W���с��w�1����5C�:J��K����������pw��b�+6�ӄ�o���p�#�ɒft���Hm%d|�4@&ti�2xm7�a�L]��_�ML��)vD
1��\d��Ȑ�=�BMѩ>Xx窉׸����4
(\0U-+)������p�Ē�@p�g�M.3�E�a�����{�wh;�:6G�xI� ��rĦI(!i��\8{WWK��T�%5��Fw��D`�x�ܯ���@$H7�AT&!�G'E�Mۏ�����"|̠��-��c�"��i�D���=ǳ�qd���dg*���8o�����ơ�ұ����26��WT�N�v��X;U��F��co�㴶2#��E���@�$�&Qn�rw��լSd���C�ua��ĝ\/S4Tds�G�bW�Y���Vї��M{)aOE}��%2Cq�ٽ�*�Ne�O�����-��\����s��=p��Uoks�`����,$�K_��)��ZI(m��/"�V._�n���Q	̉����1ݵo�*�| ���w�������b�����f&�� 0���^�1�'D!�òIq�W�_���+��CE��z�u��$�0�C��F�5�,y*L�i�]Q�9W��3;f��v.:6̊UI�����
�Y����