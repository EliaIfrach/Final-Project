��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��-�ro��i�����/L-�U��lOjj�l]I߫�p3^������_"�'j�ʬn�*W�� �a��;��}���������)t�X�|�r|�~U���;��k��2��%�`�	�c͜��d����/�OB��*$�K�[�>�)v���������~$�sF�]����ZP�6͝*����ĩ�';ɒr����YU�|��#��Yq���65��~�Mduث6z\j���4���E_w3�Cن̷����o�I��Ƃ�G���~T�VO|�θ.YW�9�����I�0�J����r�=fw 	`2K�$]�NF^-F{Ux��L.2OP&~����k2���S�BY�F���iG�H�E��+�%h�<����I�[��G/*/�F��➳��nZ�W����Y�o~r��_�$��\����f�M8D�o�OO���"��D�_U�@��MC�`��.4W��ف�O(��
��,-�h��jn<;���#��'>�鑩�!i����8�1	ZB4J�yY����p>G�����ٯ�`����?C��?��=Y%!��b�IWx+����Q�XjD�I��5��� \�u�u�@n�X�gs"ݚ�i\�X�8�xt���'� �� ��\U,��P>�Q}�������g�]�JJM,��𺪆l�
��z�G�+�QeE"�<���?�PS��"V������FSh�Q��p!�o���M|ln�P2଑��\v����7��e5h����p�C�M"�-�v��4͵ȁF[�=0�$^WHm�ضZV�#�SQ��O��xX�N������C}�4<
. ����'�L�)4��⃠iIp�9wr0�i	���{(�ĤH�:��j�pY����f�*��h�o�C���8C��,�R�����Y��//�� �s�ߚ�y`w:@�ڥ5�r�F :�Z�լ����;��$����u�K�_��B�ĺ�S[w��9��\6OU
�-໓�*��oX���M ��&	P�o�׌i�o�--^0����g�e2���د ��m|�⃩�����H��	���T�ù@_,��gx�-��[�sYa��D%"�>�G.��0y�"���(��x��E�W�^ئQW'��~�Y�V��h�P4;�w��(VY!,n[��龚>]'*�Ty�tB�+cby��	4�A� .Q9�Հ���5"HXf��f���oދ��t?�u�o�I!ZĨ�,<N>0/��4H�e9����X�C�ck�@i�L8F^�B��#@��|J�l�י�Py��D)����VV� �m��5��Y�X���
�cw���&����I���2���m��Ճ��� $(դ#���A9�&�����j�I�$}Id���lZ��ƾ#�1���%2��i�#LxQ�V�����#�J���������T7C��5��Eo1*�u0��N�6lL�d� �69���əΐ�,su�U
�xÒ#P��G͠	L�<%�V\�J�45��(������֧]��=_���]T�����@�W��tr����S�E���L�4`%9⮗Pr�ӟ?�2*������m��\P���X�$�db�mg���x��l����G���#8)����~����8dK�u�#uz=�@r��2��U�O�� ��"j�$��0F�c���G���H}�|��p{�{��ۇ6n�I��^���M���'�cލ(D���4Z���y�1�tЉ8^ێu�Ka[��fM�Y�j���#҉���'�ޢ�Hk2�,��ijdT���:�BKY���y�@X�o�d{�G�|O�j����D"z�Ǫ�$�����Ɂd{��u���K�
�[2��������Z
�ҙz~wO�:�Uӝ�`Cr��M#|B.
o���m,:�6��8�$I2�[��ll��y�Y��,|�
Z���U�5��3����i��w��Ӑ������A>\T��_�q)�,�ݒ�J㇭�ժ�P5����M��
�nW�#�_-a�)%�$���vw�9��#��<�4Ɲ�+R����������
-W��:�L���=�Rɇ9U����<�0�x!�e��@=	nF�=`�쓀,�XB��`����\�$k�j��Կ�ҳj�-QT��.2�����.�F �ɷ�?T[#B�^{Ʋ��|!Is����G��ey9��8���N�i�@�OQ�W���f�E���C�h<�4�.��B۷3����+o�drD��K�,H����J=	����/5�ƛ��ChX�0dvf��*���VnW�����!���%'�m���O�,K|���&�g����aAh7 ��e,��UX?tE3'�	J؋�`$p��)�A��]��G;�}?�{�*�~�3���^f�c����脁t\?h���b$�L��0��f:X���?	�@d��7N��#ؗ��Y^3$E৻(��]O�=�ڈ1�ͳ�k���Âq�\��	"*��W�{�?kY�����3��9G����u[#�۔u�}�;.���'��/�����",P��*XO�[	2!����&	�#�?�dD��'	�xT���)�V���b�[u��j�e���qS��(�����MOw����E���Ǳ%�����S��������P���}���~��R*�)����]aɶ��L������sEy��<�E%-0O@(��u�4uv�u>�j�7�t�)�GE��a�-(�s����W�i�`HA��o�1\ޟ"�kdQN�NH�&�Bzq�	���͉5�>�@b-� .�gJ+�!����/#h��<̟N^5�K��i�86�ߓh��}�n>I�9j7#KC����v�+�~�
�\|�*��zgШ�9�(Mԃ^8>��<C^���)���Y�Y8��:�����5B�>h^��b�0%�oM�E��Ox=!<Sǯ�%��]Ȳ<�{�9y�L����s�^���q�Ae`'t��	�NHL��~y]ng�xo�-SI�t�p~��7�I�ƲB����N��DY�=b��:�K��%�!�K����ŉX �8���*_�t2.V��$�����fա��l@�H�z�m�H�L�����{�����<gj_�1��S�SӤK�sl��+��]�41�oZ�}urW�G�2~�X!��X����g:U���H��C�/i���Rפθ�=��շ� �e0x0H�+S]��>Aj�]�_�]���F���ݤ�����V�N�3���i0"��8t(3R^�(�`��8FW��+���a�h����Pi��\j>8Q�ϒR�������Sz��T�/U���ų�����pƅ�-��PZ�7>d����.��'r�H\�<B>W�ԆM�/�^�����Nq?�*��a�R�u
���KΒ��~��
U�>������&�\EH����}QJ�q��ߩ�3�(���M{^y=n�r�C5��6x�rR�̠�d��!Z�G)hMm8Q`�q�d�F�qx�&��1�K*��n	����4/Cx	�Zu�C�6���?�#voFo@RvYB�P��Th*S�5('l�`�q���w�b�Hj;
ᄆ�^%�k��L����U�L�񍔎[�T�O�a���-�g4����M��('���+�~�R{|����rX";>z9�r�ו��Gmm_d��H����  z��~�
�f��C_��C�u=���Xr%!�%i��	\�r��+4*k^S�kpG�٫MY���L�(�I!�L��n�ꐦP0fFv�ǳ��9�0:@ M�Ě��^p�v�n�]�,�#�h�У��a��)�J\�]����Ǖ~~
?��{�3K�Lt�QR��Z:���-��Bͧ�"��m�� e�*M v�uљ}tؘ�/_��,�T��Uy�A�j�ބP�S�2!�V�MWR��4Bv�c�:V��kݞ%{�Y�>n0(���s��i3�pb�Q{�l 1�S��|y��r�������1�3(C`� �;	e�O�B�����N��f�w�����k�7_3�&����Sk�B�F�uc��M�#i7y�yL�dn}n_��&c]���!~�Pr��jU#i������a�������~�F�E�U����o�G�e肚�aMKs��H�@×E��-�a��`�<��AI���Uy̍P)�!�t���D���ҵ=^
ϼ�P���T!Z�������_��I��(��kؿH��������mş!�)~��p���^]�������,���S���/O[y�����&4m�k�j�*C�G�yKn�j���z:�51����'B��ߪ��B[�Ļ����/��)���xQ����dr
.y�ݼ����*9�`<=g>���^��U& 7WL�)��JT�W����n��<�fVxQ���!�����#���0{�֭�5tA��y�:�J���5HE�yv�ײ���D�ueZ�r)U�c�B%6��&:*��#nWt:߀���L"��Z�a�/�f�%>�6t��N�mK���G�Y�xyWL�ܓ� �A�9�sg~�4����G��x�pC�BW�gm��,/&���(c�ЌM��:�>��X��H7
77A$#�:uIH
�m7�R�[���L��`�_��hj�����XQ�L�2#N�0��a�{�VӀ�X�]ء��E04�n,4�=�E~q�E���P���%���5A�:����i������2[����q*{�!�v0ii'������Z�~����4!L���~��M.b�)IƦ�*�4���~�t��W��`zq�N�m�+e��Jtc�8��zgϓ�m�)��V�&����I� ��|�1M����:�$�OdGVL ��2�����C�A��
�r#G_h:�
XSx��j(R���	�&���@v�ZW�^��<:�2A)����,��S;u�����|���K-jH���6��ެ��z`�>Ŀ�������.l�A��6}�'�bW�~�f�B%KyĻؓ�[J^���G�R�[�&���vS}A�..��Anh��~��v؎�2����8F�c�J���Dv�^�H���� ��bmi����	5��3��b�������o���z;A#ئ�i��~������v@a��o�%LE@z��ʎ�Tq׃���,·#��N51 8�6�(����.����'����$e�K��F=�J���+��2��{��2��N�#�6/���~Y������_@u��1��.��Ė4 �E�����0�0|���a��l��²�Tdge�JՆ��t�PH�!�`b雚qϷ��Ƭ`�9e�Q�PR���:X����Cpi{����C�H$����r�O��C�z&c,l#�fF�?�uR�_��U�nl��2: �8�+R���	(�b/��Q�Ā��^=
��Q2�KW�X�&��a!���	�6�k����MoTۼ�,\���H;���^�5��4��@'�
��Y��F��^�I�Y�-�Β��L	��ycl�B��nz::������L�U�.qtS�a�vLq�� �U�M̂��f�%�3}�����k������9�8���l�#���#���A!��"ukX�=Ӌ�Tn�鸞�#Dh$��N����Ћ6�sH��P�m�ghNV�l�C��6Υ�H3*��
@�8\�\=��Ą0��H+����^�>�~y�]=��ݐ[����<!�1�H�Rw��c���>�a\C��z܌��RRSc���G�z�5j$)/���Ψ4�ƞ+Ҁ���!ضW#�T�������u����4b�\�٘<%�>'���ᙴ�þ|��\:�l?�6��>вz����F:�|�(Fs�snM��`[j���J�j��*?c�����Ǫ���WPW?�z�Yw'�ݳ�	�����h�#�����Ĺ��[���Yun�YA�?�F�����p�O���ϓIG+���L/�#�m�{
�~�3�}�-n�3�I����xnH�ض�~��N��Z>F7Ԅ
�������^fC�;������%ύ��yK��>�U�-�}�������$\�r�lt,�j����mAx^f�~'��Ӝcm/��C�� �����/?F����I�S����5돩.���s�DbBt�I���ԝar
�́����:�g���l������"�-v{nl���%�Ҧ-��)�ߝ2�r5�5�/�C*ف��4c���9��NVq_ť��M��ݾ�iʤ$ù���K E&\t � �dYx��m\�����+��:pLT	��M fm,��џ�T~f֑{�)�;_�� f�ތ�1���ݧXkhӽS��"�vN���I(�?��:�����bA� *=NW��#���f�m
��o��2>*�iY'ĽGx��O��n2�^����Zg��ld��݅��,C��3��L�$t�E��
�%Ko��a�M�h�g~�Lk���I�5�W�ݰz:���:��TK�P�rR���})|{e�o��z+yyV�=����_� ��U��w|��Gz|�>���rI>˦ o�.�d�����v$��m�ѷF���K�~����sq�x�����g�戮lţ����jz�/�	ߢa�:@�]no���>E)���A<W���KH�n l��Y!r�i6� Y#����*�F||ޭ?�7������vfK#��\��X}O�eꭘ��Y�^g��.�[�:$S��\�KV�U4������I�&TP&0i��K�#:O���:��Z�56�o�e>�I���cyI띟��
�}�~�����ƕמE �J�z��,��n���Kj\8 ����6�߻�ɞX�9b�Z�ߗƀ�%/��o����UHr
����L����?]��^Ƚ����8�g]a�i�-��r>���O�}�(�|�F�V����d����zRH~�|��	��\�5� ���~ل�+���c]ID�3j�����U��Y��<���}�mE���8�fR2�N���1�@�?�쵮����k�Ql�P{m��$>�<��B�j�\'�+�����W�X���p6���=�˖��
4�s[�����q�����=Z@�[Z�VmY9}�\���H��m"��V{�e>�c�V�:|��J�7��э�����Y��y��\�i�
yx 6n�|�B������zpO�3����<�i���y(4G>%{`�v�t3<��.n��q��R�"p�x�RbǇ*�¡'�J�!L�+��58���}�%j���9�L���Q�'��{�: 	��1<�k��Ti��a����R��Ky����b���-��������_��Sg����B1�I�_��E'	byƦis�ͧ��Z ��qq<?�_jDeⰤ6r����M��?2=?F�={(kuq�<��� Q�z!�%M'�_��z����i��:7�w▂���U���S�9���|�[��4�{#�V�p9�9(�[��؀[��<MF��<��K;��(	������2k}�;lV6�ޜ�`���)3O�ޯ~�m�*��cx+U3���"_E��^���*ά���5,^���TB��l��Y����A��(k"q����Ar�)�`��pD"�#�֭w�����F��H�"g@$�x%�y Jx�Ηr�y�^)h�h��V6�SNd�2�M��0O"z�;"`�ƫ3ӌU&0�RxF���qHh�:UCFn��ٽ�a���SdӍ����¹�8j�x�������3?�4&?�@{�Zl��-���,��=_S"9>����U��%L��"~�y1�sn�Q�ف@�P��Sr�d~L՟G�+)�|��IO.��\|31
~�F;�'yW���{��Q�w��P1�ȵ���BH����)~�f9��r�,�<�E"ʹ��*�k�?�U �Pfڽ&ON�%����v;ڔ8�l����v0�ķ~��3���d>%�u���]�� `%�Y��ﺺ��(م��S_�z:��������Ȥ�D��;�\�� n�fs�4|O�Nm��r,�Kg��p�X����X�����P���ͼU���ҿ������L�m�fS���ŗ��c��k��݃@�nj�~���QT�[DO-#}����Q��FvKK�k�>����N��S-[	���'�Zycy(�����'gf�D��Yx�E]�e�X֝'�׊FE��<#�mr�9�L%؇�(bb����M�u����/��6�V��I�[�ϒ�UY�j�4^�l�M3�9�S��0:�9Mu��8��=m?J�k���=�.�(򉴖�A^:�����kiA�����3Voj4��׎)��!��J���|[�IC)$���lF8P�v���b���I��Nb��������)+�,F�;DR<!��U��2��~�7
��̴g� Ӭq�v�,I@�lS�I)^*p��
M��ߔ��˸�1}p�����II�!���?,�9�V+������Oߖ�+�{��0�ŷ��skEh�.1��6�b� ϭ�SI1f*�&���z�ۍ
k܊����A�"����vA�P8�9�m�{@����l;�c��<7��HV��ۭ7�(��z7J¾��_��CQ�4@cW�$��$V��}Y��'q Y�VFk�H�q=��P�u�vx��ru���-8,g�WVS{�^��R��m�ט<�M-�fF��	�z1Q	��9(�t����8p�R08Lg�#�p���O^��7;�:T��,I�%"~����@�n��ɀ*�*Dё�gp��@x]Y�Ǥ����t����������B���BӜ\���%����ya��6��\��Z��㱫���7*�m�U���!b��?�S�,��j��>�=��dY.jh�x���;��T� א*Fx�EvU���ǚ!�P[�?ٙ&r��񥌝G)]c��W~g�����i��C��f�4Ȏ���9�\��:�Q���[���*IVz��-�q ��4�ib��'�P^z��z��.x�
�6#��WH/����9�:��{`�;S�.=���H�����W��X�)a��� [�~�/ӣ�B=i=��µ3���á��&�TZ]AT>�d1h��j� �v53a��b�^��s��n��B�&"�����ڐ��L�C J�T���3Sx�i���^�s��]=�Q�g��gҙG�`3'��إ_�G�y�wc�=g`҇b�c�䱫�����nߺփ����DJ%��i�9�j=B2X�z4���"G:���ZԮ���Q=���_oW-�sy���ٯ��,��ޞ9�@�>�U���M�Zо_ �3�=�\�`��6Ot�H�	��Fm\�ȋ�u��5����m�'��Ӧs��t,��%{��X9/n'�tIC�Ffy�̏E��"��U�P��1H�U]���s�>���SP��v�����n*�-�A���ŬY��Bm]nضS�dS���L4,� ��ּx�Q,|��rEZ����� 6��ߋ�g����ي����5�3���fai�����j2�px͊���8B�����52�3��/�>�&�tX�ǈ�����s.���M�X��\(�[�4h�f]�ɟJMw������T�ET���qu�$��	�t}�ȵN�����*�`
qL�
��|v@�/$Zu��C'�@���=�M�>c*ȉ���XS�]��q	f�R��'�L<d{#,�@������'"�_��4+�=�(�yT����y�% a���^g�njN%���߁�jŌ����MV�v�fr���@���lh�4��@���?썹��`iUsu�o�ڏb�ntn�wP�'ؒ����K�wz�y _�jL�$g���������'�/��}S�8���F��:���>!�hG,��hZedӃ:
7̤��?�,���L��%*��S��Ǎ4�E�HHJU0g�>(�`|�M����t�jC�5�~me��F�p��8�g�/Dt;�|��th^kS+���^���1��6s7��0a>zaʕ�K�hx��+�`nQ&Eb�]��QfN>
�߻�q��j�����r\#<�=�"=�XV(w@[� �����"����6 ~@?CV�@2s��G)�Mz���*�!��C�!��p@�逨5g��<;�>���x�'T�~?���~\�P)�Y��N�����-�L	��}���6�?AG����De�Qح�� Y�p3�����6N<�p�C���'�`=���0�����c�(YY�$��k�60~�D~$j����6:�jPQ�;L��q�Ǳމ���/�)r� �\�?���e�F.b��]0��N74��yc,��#����(�>����}F�|z��4bp�RGv�iHj���[S�V	��L���앍w�E���yrb�U�TK�#+v�������T�bU�^�Ƹ��,��xLQDT����w�����*��,s�{={��/�Ba)Y=�r��(�g��$n���׼qu�	�[L��(��ּii�k<l)K��,賏/t��􏿈�c"O��-Y|�����Ι�=��IS᙭��b(�~U#V�Cf�dH��b\ΘG2�lK�>#Ҧ�a��0�3ԣ\�Al-���z���t�;_�t�����h�I�r��keG �Q��9�@9E�Y�aw�Qإ0�kE6�qY_�>([ڙ�O�]8�Ð�j�M�H��W������:+`#��c���=$'��a��F���ł��7f	W�\K�1qK���|���S6�dh�'qW�"�2����d*QF%>`��;�7%��W������V ���_GC<��*oF�+��O[����H�q��-�<l+07��-]NWa�I7j�{W�d'�8
X��&ɗ�.4�K&`�9�u푰��T>�Ӡ4D0i��W�;bԠ=���&Ȗ@�fߎ�H�����z'��a���2�H۔iG�,mo�*=��rad��\�n�S#��-bF>���J��o��=�+�@\�^�._q���W��L���劆�Q�އȈR;�}Y�g<E��]��hl�f�i	,&�RZ���l�|a�W<1�V�3jſa;�#�)Pf�[�$�[�$g���ʫG�dd#zov5abwίރ����\���|��E[F�WKh�0[�uH�lJ�C�[=>ZH�`�GvD;���s/���6^��4xH5{�����$�?�C���#�(Z���cF�K<+Г܊���hValv���Vq�A҆�;���z=x[]���g���9����ŏe373��`ɔ�ݶ��a�|��sÔ��G}��V���������>��E}�&j8�YQ���e�G�{�7�	��Z�@���Z�д��{�`���#��*�y����j��X_l�=G\m=��q<��G����A��컚MW�l��o�Պ��[���Of;��K��N��f>EYfq�D�6�!��{ef�k�
�1�9�����΃��Y��N�7�7�ͦ*f��KStzu���rc>�.�[h;��{���+
k����γbPӃ����Nާ_��N1���ʇj������@ֳ �͒�s+�<���]��#n�(�Ҏ)��BHz'C\@���e[_�!0�ީ
�Q�y�= ���n~�����*-HUK;���^�*��Q�kb�F,��o��:)S,��Z�V��ܪS�(�Q~�ޒ��@�A/���J����a8:�44Q��ʗ��-X��!s�Ln�y��x����!j��mA��!��=�;��:US���h4����_j���1ޓ�*E��-䟍��JY@��mǀ%/5��_��OL�PO����x��٥@+�'�5�E	v��J����g@μ��7/��s�^�Ae�s�J�Hf��ApTv�3`�����{��Q�$�p�,r�Ʊ�*���b�{��s���^lP��S{�a;��h��OD9��.�J�S��G,U��p��a���E�a~��Ic"�t�S�wC��zU�ؙ�08�٭��T(=������FĞL(�TbJy�\\-���j�Y녍o[6*-@�>eZ�Kɧx���ް�HLz�H_�VK��O�K��H�zv�K��F��[&�̫'�ǲ��V-ib])u�O��
���s�� "�I��)��`��r��b}ɪ�Q�\r��K-% a�t��ѤKJ<
4jp��� ����5���(��B�	��kt��<����e�4�����c�j<d�!25�b3���ho�C>1���&8�y1MM�ƟS��罱�C��S�ӧ�5Bj�0vs��t�j���w���(��d-4�i�,&o�-:�ug� d�oa��T�{�J
|�N���Ka]��M$��9���y�0�U�{�	��`�/��������\��j3�B.�@������St�� �M����k�u�����|�D�������:�B���A\�戝�:�r�����R�g�*m�3�8�$�J� \�{`Z}m�jG�y�bʘ�ͨ�y�YBG���!��qY��끺�
FRd��m"�s��AgTY5uKTL�!�J�%�����Z�'�PA���"�X</m�p�~m��l� M����*��
u!�)=\�2',lwH�i���M������w]m�=W	���n��D�;<�^H��
�(�0Tگ{Fdt6ܭ���o\��A=Ʀ~4'(�Ш�afKz����$��FqX�c����x"�:�O	�H���[nR�-��X�֖w-�m���c�9���g0O1�&��c�ɕX��w%|f�{ϧl@��/ ���]������O�@�2�Ǯ��t�]e�cR?��Rx-��]���ԫ�1�_�	wME��h���8'qɟ��5���s�Q��!؀��#�֜
����ى�q[I6�|�� �1���P��F1��K�����~b�C7�4���1�rv��]�H�i�Ϻ^�eT�b��������19N'��Aڰ�,�2�TM�iJ�ē�~�2fnV�'�&����5g{�AF=4|}�,j��M T1�އ��by�/I�A"8.��zPd����: ��sô�~��&�ԧ8�v���vk���"�����9)��&�^����G5��V$�瘃:U����U�"��*8��ˆ51F�3��Q����EM�M*��g�8\3`�a����7�6�n��/1p��w�6|*��A���G�ԉML �r�:�L�+<��h��М��5���'��z�}<����c�K��_�~��aJ�(Z��#�:��>m`C����@�"'���ay�3��1�U�3��3ށ&����{7�Pl����r?Ѩ�zؚ�\CND�sk&�Q��ne�0�ʨf�3�������O�$ᬬe����"}>�+��������O�R�1��5�e����w��;�CE��l��%�
b&j�G�~vl��$t_YCE�н.�=��8��.A��uq�̋"��1�����*[�P�$�m���rV�&tZRA��ܢ����{d��vn��"�g��EIE�ַQ�q�ѕh=<���+�b���G'N�;y��:%v���	�+�GY�.U�$Vt�������9zr�MYe��y���,�?�Z'���}���?JI��z�~O����hn	���G�P7ڰ�YS���1I.�Eu�2�r��)�%?�xA�?MG��v���4���\	�|����0�xį�I�5�| �`	��K��ql�~Q�W��8�.ϧ��֒h}}�_网�Rq���|w�q)#��'�m��Ǜ>�w=+d�\L7Aй/�7�t�u��E�yi��KЕ�����V����s@���Q۹c��k��<�b�xhu������Կ��o�>gJs� k���[�@�QC.��+6b�z�M%���H�:��oױɤᎺ �C	"�<ht�.:#�]�ȓ|���H�o�<eRU.݇��\<�huf�=Q����<J#�c��Z���8F��@�v�\}U!J��}|8�?�� 0���6fM")&&)�N�A#m��r�3d%��L�$�GY:]�۾	E���MbQ�]�H}@*�gY�����E_����~�\u��|L���R-:��WB��74&} ��Y^V�I:��b�A�a�B��-h�1MWns)���)��c����z��+̉��[D��P�[��\va�i��4pb?$���d;Ŷ�{u�~�q�����J �`���c]6G�W\5���a6ܥ�]�� 'c �����C��
܇n����o�E'��Y�g�4��A��|}�Zv{p�|��ק�Z�/���p�9f	n�y=��j��x�c[���M�,�=��	!�Dǋ����G��%E�3$@L�	X-��z��殍[�(����3Smd���%�}n��SF��.f
����i������	��
�\�dFʘŸM�	%�YE�%��L�ǿ�6 �ݜ�I^�N\|�n$�k��;�o*�)x�8G�ݫ�U��>�S��>��W$��p0�/���G���g+}���X�+�3���uZ�q1O���ٸ��M��À�zT ��=BΚ��_l�=�g��������
�Ҟc��L�b�qU��7K���;�`z(u'a>Hbl�)QA���[�4���n��mi�	6�+V^ؠ"č� �=��n��_��#�T��Q$.�0�IXǇw��P��P�Ķ������|񌭄���	}������2�13��jR�ܵe�" �/�r����%Q�Y^=����Xdw(�. �Ɛg%B�vX�33r�z1�O�n�ld~� L�C%�ET?��튺o��y�6��߸A]6�}�ƿ(f!or��<Y�{Ÿ��Ep���Љ|G# ��v>��ȫ�f�����z׀��Dn��L��%[M�\�O�2+�E�����*n�
�(��\�\�Z�cbB˶؝4B�[s�.WQ�_�X�.���D$6!���k��4e��6Mf���[�]b���w$��oJ���AU����jsE� �+hctxv����(PO.��'X�=߶"��J��ݦz�҄�&:��3~��RR�Bq���]��`ǭw\Ҋ�b5|w��8�����+paS������W���E�4�.zk�k ��+�1].����1�#���v7�fS'L+mG��R�dU�
�7��N�K�H��|���6���������{D��3nRB�(��A�e�����U!,Q�� c㉴;�RH����7�n?� 10FEӦ����5�ʟ�
���J���(�f�[F6�S�>�������j͢���1��gػR?�N�jQy�_��U�g�U��X��X����G�`�z�.e\�g`��h6m�Eeo.m6���!IN=C9�1$c˛�Wp�h�>��\jL�|  ��fT\�,d���� ��A��]Rr���R0�G�G�$ਲo��m	�Q��\^4�I�e�~�/w��>U�!�agu�����?ȊO�z��U�Al��k8N�+�QSb���,�����E��D����|~�������`�\6U� �j�c#���]G���P�-g|��%h��R �n���!�����a�2�]�����4�tw�V�*���;l>VZҘM�⪀m�C�c��Zѕ����V"y�2:1_�Q�Ҁ�k�J)R~3 A�Z�W&E��$*�R����A6"�*I�F�pi���?�	��L�q��|��`�Ez�F'z:p�w��S��RU��FX�YKP٪�ˌ�� j�� 4ei���fi�<��E�Hy�҂�FD�1��њN/���3W_#�SzJ�[0��On��>�x���S��A�q�l�K3�V����9�9�EqƝ�]�򋴪w�nS�˔ ��C�v۵Z���u�.%��LF[���L�M# v!�y?Us�rX"�.݈q<{���B~�-R��j�ˑ��p
U�>
)<�KםR�at���{�o@�K(_(i��
��X��;A1�0��7{�7*��_�	%�sjn3��olh����!s�c󁶏�E�7�w'+΍��f�~u�C��}�m2�:0!ޱ}\Z�%ո')�ٞ����7�]�`�4�k]��� �[
k�R����S�S��RjL]�M�y���u�H�-�ykA� ���4G��S'�g�ssR*pģ@ag2O+����T$ [\s���+vO`��
�2�,�ͤ!&�v?��]j�Q;8�>�ƫ���v��@L��Q��I�sʐ7#a�V�OɺJ<]!+�� �ExDJ"1LWkϔ�V�<����8��A	�	�t5����� R�������G'�pf���L>�x�4N�</�<���@��G��n�o�
+�1WK Xl���}`�S�cIfKp�R��N�]�^�?H�?Y����{���׈Z-f�����8-�b2ha;UNH"nk��dH�;��Q�ԧ�	�y��*F����VP!Z���RK[\Gw7]2�k�*��.�N���Z�2]j��#��Q0*𴊫�9	(d�w�_<1�t6}�G�k���!�#?��	 (���l�v*Ӣ��g���&6���If��k ���vY.2�|�Wa�G��M�����"��ٳqsӝ�M�a�PLL*OJ�j��!�TY 
c_�3�]�Fb/�e^�7!�Q���:�m���J�4�$� j� ��T���Pv�]�4��9��6x�U���\M��~�BK��L}����Fp**ܝ�6���}�Z�ܘN�7�FeĸP�61N����\RP#�6���'{�lE��+M+�<vZ|UW�f�+ѵ%~c5�O������}і�m%|X�R^���X����g7?�P���!�Y�Dk�~<3�O���v������,�;v&w~�5��M��^U�w%H����=�O�(�].�)`>Zi.*���D9;rM�(�wl�N�'>����C�3k"{,$&�T�������YC'�*��R��uN�$Б�t�;%@�6�"�5�xa�r�`,(u��l�� �vM��K{��y��h�Q:YH6ۈW�(w�m��K@K���\v4�n���v �T���4�+��vRC3�7d)���;,>��X�4q���<�ί��O�G�ct�z��}�yL��}��=1s�����LW8.a}�З�MK����؂�D�-�1&�H���H� �)|4���p����"@m��*@V��V�c�i/O��;;:|@2젖��̏5�4_c�^ɻb�?���6��w�cX=s#ӱ�cj�$t�q0����3�Y6M�X��2���h5z��ߞ�CV���&����a�S>���/?Y���˙��b2����E���y�@�Qj:�։{�?��xTX3�=�qG�/cz>U�)?���cz����E�V1(%��a�?�Jw��ȏ5�9�ܒ�T�em
4���Y��L�Vzd�D-��9Y`L���$S��4.iXO�
����#�����[鑌s\�-��:�w�:��8]�S� F-�Z��PrҌ��#�H�
��n��nW���%��vP��7��`a;˶�$M�'>� ����ώ,�p�U����jcm�>j<��Bm��?	�\��?0�R��/��ns�%�M#9�n�NQ0�9�Z���ӆ�v��[��!��`-T���ON3C�z��@Y*��>E�Ve�]��t'��E�zJ��Hq��eN٧D>Ұv��_՜�A�7������	�(+oГ�0���`��$�8#.�?�?3�NTZ�/�H�R���d\_7#�6Eϩ2��j�}����+a͙`���͝�
��+����`�EFMr6���1 �L�3�&y�ʼW���D��KPG��(�7\�;�P+�bW+��+h&٧DELt�Ko3�lZ��)�Hz�����9��W�]�=A�5����6��tH5�-A�G �ƶU��y�d�~?�ɺ���ڠ�0btd��$�շ��l�6��#�{�tA;Q�pX�Qa � Gu˷ڧ�4��ժF�&�j�i��cl��S�e��oTht�s��S�q��מ�D�V�
*�V|�JP���"(�:�ѐ��I/W�S�1b��(q�HV�?�NkSj_��ܦ�K���l�4b`�bN�E���Qe����JG1mCɊ�Mj��7�m�����+a�ข }uZ�2Ô�#7��ݧ�y�b
��sgI��y��X��"�� �_��/7�0#�v�l.�i?m&��<TH��B7�%�����k3AB�X�����W�Vf�6+��bc1��T����B��d�V���]uc�mv�2=7�.�O!������%H��A���)����l1gت�4�HQ�0�3[s፟�����7�	DT��W� ҥ��(NY��n m���MC�c�-�#KnD$�Te���R��0^/y��������	���[*�꼝~����zG�G�2C�Q.���On{�3��jZ,|��-i�����y1$��bS�:@�HɅ�v���R�q�]j�`5�;��Ob'�v��7t�R����D$+qλ� ��S�1�O��=�_6��[�Q
7UT�^�����aL��`s6��걂�vwυK6�ч��\����{9E�,����� p O�Q�A����5b6`_�0ŧ�P�X�#��ey)�N1%��)�a�e�Mh�{6�äk@&��RR�g�oa|�W
v�!�q��4ġ��۷��E��������ȩ&���.�6�5qjJFD����R
c���
��I5�G�~`R����W�:B8�T�껊ӏ?�dЄ��;0	���N��Tn�fp>���M��g��41�R��Ư�5J�	� �x�q�<s#0'����_t3�7�c�Ot�|�8![��-�>�ag���Z���!�/:����i[��.�bz�0���@z�d��WX�l�{�/\?��y� �;W�E3(�/��:���V�d�6
���n�YJ�pb<�lI��X�]*���@�|�F<�����κ��Z(Si���~�m�4�(�u�̣�v%!+���0s�|�:@u]��Ʌ 筀'ą��Z�y%�)�/a#����M���}��8O�eu&���-6<\�HSi٢�nL���&�q�1���B���Tp��a���$�Q��y疲H�+A�7�AVΙ@���'�I�5H��"-�5�&)k�c��?�Rv��#�s#]vᒧA�%i�	��V��2�����g���4s�̬����W�[�.�,���x�쵝aqB���֛��%��������3'cQ�^U\$��w U`m��V-e1A��`���ɦ����A��4���u��g��-�ҏ��
�m�o<��A�_*�03�C��V\PC��o���L�"��`�&�1d=�v���{��vO�R������)e�������L�Lir�RK��<�f���}��^�z��>`)�3.h_�V=�|k	(���{%��-[�R�n���?�y�E�� �>o��/{�(,.>�C������(��B��dBLk�(��N`Da�,��a�� ��=<t�[���v��S��)(�"u�L���lU�<��m�g���g�
SH������&�o�իw;��W,�? �)�������7��5aہ5�� +Bx�*AL@��ގ�"H��OF{��֕�,&��ż����
b��6d��$��!]�����lTZ�VG���q�sQ7��c�s٩�m�a��f��q=����ȑ��CL[N��JD�uw�
c�ֵ�UI��*�g�	����b㱶c�y�WT� �k�)��	�)��r�FTe'է��N ,LC�t��y��xȬ#GJ5�d�8]�SEO��K��n�\~��xi�O%6G@�^&Ň`{`\N��wДy%��K��%����v�h�۸ Xd�yY�R�ʧ��U��0B�bH�Uw��aF]ͩC�+���)W-d5V��f���Z��'9ܩV�~*GyG�I����{�5۪	�ߪ9�:D�%�-��:"��4�s��z��VJ(�^����f����8�d��ɷdJ�L8*¶�L�7�v+�A�U��nm1|���.��\�E��)
�q�����q�:�����.��h}���'`%���8^�,YAψO��'�eMcG�U�5��iR�n��t����Վ
�	��xf��i�_��Ɲ㗢>�|/���_h�:;tv�<��(:�v��R��,���8k�>&�a�ݚ2"?]�Т�ĊZ�mAwgܺY�j7K���1�]J��W�j�K�h��Y�\�"�Dn��0�5E�`3�
�BVQ��e,�,���e�]ķ�q�8�1� ��C��f��crnAC��t�~n����:���X>4�[whZ�D�ȸ��*��³w3(�P�Z8�FF���U�F������ ]�#�ͨ~Y�^��ޱ�]Ow�}N�Kе���p$���t�P�ؼŶ��Pk�Fv����z��f������<ײp$���t�n����X;��?�˓�ٵ^y[�{�ye����zQ�N��#���ݣ�ʴ��m�A�߼t�S���4U$g�&!-��C���aE$��4�- ����N}$�T�i�ztt1����-�riM�ܫ�pڙѝ.���L!�.����d4>Z��[����I�eeX�(���K��n��*0�!Ye��R��[�vBk�+����@�����e�Q�)��`'.o��ԝ�ە��w,�0�ѫFG�g�"�5�5�r��^���N���޲�Pdo���t���K\�p��>+_������sW_9>�`r���t��a�1z�],�=I3��a�wq0�1��C>i����� �q�\�:gb)��c��ly��<@2*j����t��
ڞ�)J��xT�����$wTg��Q<��IΆ����ۻ��c�KJG�*�m������n��+; �� tq��S)w����������'f@�X`)W��g<�hwM���\���{�@����6�u��:\X�����ɝ9"�q������'�3A�y54���A�!���3��w)�����f��u�q�/�>�P:��Q;���F�=��/z+�e���ܷ��3��T�*��W�S��god|9Ž�G�����6��$���dd��L������t�S��EP$Oz6FS+��0�݉"��%�>�]�~C,I�v�Z����{��!�(WO�
�悧r}M�G(����ج��]��e�Ofzl*$�4��-;����ٚѠ�+�Q��,
��#+�| g&����Ay�Q�5�b��1��ܦ�^cLO�[�w�y7�_��y墽��|^��`�I��x����`<����,-[E���pc8}�(��)x�y;���{=d3-e#tnq��X������p���.r�3Z��� \���y
�fگg�M�_�g��Q@1��5��,�7�/+�S�ܟc����=b:s;���X*���@��a05wj�}!��b��K�vrs������L� m�;�� �9�â<�$C�H���1m4-]>zCiנ��Q}�\vx�&���(���t'o�}P��P�9��&�p��C{���k��;&��A�8��;:9�,^�d��]��N4im��I���.���ѻ3��`�����U_9�t絥]��3��Fl+ �s-��	�Ehu�����A����ԏ]�2����3�krQ��>�O�W���ܕ��������<�c���r�� ��DRV��"&�O�)�m�-��L������s���S$/z�����I&T�r����A|�\ҒϨ�ρ��B�qME�Pb����2 z'�������e������NA9���?�*�X�v=Y�L����ƃ�\o���e�W��;ĳ���.�����W�6%g���)����&��>5��
�CM08ψD�g��n����������fj�m[�TD��Q��Sp�搠@$�?@�:UeK�z9;ON���!�'k��Q��:"w��N�PL�v�(-�Qw�(~]���0~�(��
�5��{#E���n���y��	a�zJ�+�==�qo1�D����%"5��b���'? F���HC���Q�٦��)M����JW�Zôv��J�B�i�%�5\� �ծ�W�w� _u;>P����<�/:��o#�`����[������}����o�s9�6N&~9�������Sa�v�'L������� �C���I����@�J�0�;��4"�yh��,�3|�h�B5;C���tz��I�y�>Z��C���a�ۍ/7{pfw�����'Ꭺ����]_΀�@E���>����j��G��9<W�+"jrBo"mI��y��?=�]!bQo�^l�ym�"A5�Ģ��Lx��؏"�m�
Viӯ���K�(?��ד�R�Ī��B5[PU�Ɖ�°�e��0�y�$�����m����T��6��2�N=8��&������ǒ�fpܺ�X��_���B�����i�"�?��M�-e�*@��q<.ҩ��z�m}u@���T��ʮ�����	�34j|\�ɑz	i�3��H���κh��?p�$�ޯ�*��7Jz��@P��U�������To)��h�S7�$�X>���aeU:-��S�@W��C*�:��T(�éG�/͏�5؋���U͗�$8��CC�-� �1G��D��'���o5!�9��4(s׉3x);`�c��݉5��}�Ԭ�!<0�HK�~Ȍz���'Z N�p����Z�[-���X���Rz ����t
@�®�Lƈ�>k͎:MUh���|��w�x�N-&�a[f�hxtp��(�`��If
��#����rt&[{:0J�
B�FBBH�k�X��UIiw�*n�o��li����O'�d΅�iTgT���xe<�""��2����d9�_���Cߕ�����U۾�?�<�X?s[����{��@���TYJ0+���M�ah�BI��]��y�T�t+Je��;����$�\��<M*�eQJ�����dc�����h���5_3\�����Q�{ֽ���SM���Փ!��AE�K�ʌ5�1O�6��B��t��"6�R�Ob,j�O���d�e)�	��������p+��j ��;rG�Ez:��N&?�nF�HS�@Ď�K��8�����6���C|���8�!�����L3�B)덋��3�\���5�tj�qv�����쭺,��4�>N��k:�똦���ݝ٪緬�F�a�{���H�x/A�[`�|1�Iku�]�b��#5l�n͢�#g��Z�Uk�W.y�	͐�+�Z�~S �Va�X_�����ݢt]�,�73��dd���2���\�El�9��,$��xA�F���qn�#���{A��>҅���ӿN,��,�s�G���@~��;^��d2�~�/r����w�f���6����3C4��!|n�a�2�H�3k��D�M��	`H�d!�/�4pjP�ZR�)� ��@5�3(�>���i{4�H�H��D,q�(z<��v���<���c���F�6C:~|����FP���j\�b^&cpIPox�;�!��#�+���Y��rƹ�L�k�&�;.8)�W@�a]z!��f�{���[��}m�duǺ�>�/Ҡ��yQ7�Hϣ�����S��L�`�jZU�-�������5�������(Ұ*�9ט8�9�6WH�:X��lFӨ�֠F��QH�a�7��qUS���~�DJ3��Ga[���}�g�������ϓS��^Y>��"�ଐ���º��� �O��%�K�r4V�"Fz{9��������e8G��>�s�yI�����2��ү��DR[fe[��P��jK��k?������k<�{�;lq�*=��$�ק������-�*;d==l"v����$ɿ��#$_�g��P���j�~<3 �(d��-I��e�}�M\ht���L&�@�����ٿ��>|SlMC����=ƿ���.�[|1����"4�AϏuFj.�����:%�P�h�*�~p.�{"9�*x���ݍ+��e}��I��L�8�yﲞс
���R�n��c�݊����
!d��cGlZ���Zk�r��<�t�^���Trﻺ,;Ďm�1$Ws��+w㛽A�W�g�y�ᓑ��1Iݾk��)�h9*�r��-�/�&$#�*�FzЖ������`g~gu t�"�ﱿ�ݦ4� �%F����%�)�4O�LR�.�G�q�5	�GBV>kl�f��4�Z�=�}�Պ�я��(�핥�C#~���c�eU�0p�9i���{SM�
����inV�]̯S�-N�Y���V���H#���̢�ch�f&���|���4������\E�fF�����z����mX���GV�����FeP���� VN��I�w�p�"ȸ��^&��j��!���b&4�)��ő���K�������c#|��Z�a=�W�Oy>٩sz3�?
#�s0� �C���7s��%g�P3K�S�l�!��S�Y���˔Je8/�Q��� ��h`"��m�nWelb�HR��Ж�^ݖ�b� `x�S�(UĦ�MRψdax�0�jʖ
i���8��qsJ�XVϺ��8��Nzw���ri���w�I���kRfj���\~�3���l���׹.RM�I�07�U+qO]�w��˵\���iq���M�����!��z��/�,���Z"N�	���4\6��!V�T���Ã};h�W�+�$s;H��q��e�a���_� y	C�4x#�� ��9B�L��@z��{*Ǵ?�QP� s�]BR��Ȯ��`���N�Aa{x�C����� U��$A:_MbՂp��^E�I���\�)�����Wɹ��8=iy���,gM��?ψ���G�5?��j���~�5U�{V���>��U38o�dt��GŚe��N&��C�h���mD���{�r*?a��\��#��\��b�
�rF�K!�w�*X��GI�zP����ҪV��7��y��o�%�g����n*��F`/���@Yf�9��T\�9L��v䲉o���Иw$4��}g$ܭ��#F�rhM}����jl���Ԉ�L�n�{[[E^��T]ҧ\��]rD�YMK3�{j{l�;�#|œ+��8*�ʋ�x�\%>�[��پ����ӹt�/�o?������5.�!�y�P1b5��J�
�5^�w���~UJl4x!��N%[�:�*�a��j�z!^4Y�'�{�p�8����;��������	Lz�m��"�.gP`x�)�������ˊcEqJyޮ��o��nS|�p����M�L]����|��2���|��^�Pп��`�;�Y[��.�˂]6�e�8�b�{�LT��d�����k�V]���>��\���]��vn u,�GXn݇2X'�%��x| V�~��V�C��&��8�����4�6̚��Ԣ��f�b�	�`)��xy�)�X�ۉo�W�1@�@~_/�������AH$���1�v?L�u��u��#^��6!��#�Z�����1[p��~��C	^'S�����7d��ҵ�%_P`�8��'���$
��g������Ra�f���h����-:)�t�1O޶���&x<�l�9��N�-P�!�[4�t,�\���}�W�DI:1�`���c�R�o��%��ߪYEE�{LK̽[���y��F=��guҹ���ȓ�HV��ҟ��h��S���Ti�}L�5߈C"�	˪�%r�p�U.������� ���?^Ƴ���#��aA�[�vs��$�����="mm	����ɻ��W*��C���`�:�}e4�i�e���;�$��X _Նx�_�d������d�ƸA">�Ȫ�8*y	�F�����������/CУ{�g��,��ԩ�#j�ھ+��c�iP�c�t�T*aBr���d��oѷ�7"���$��O��2�0�����OX,6�$0)��de@ű��S�e�R�덭_G�W/tsz.�	a`@0���40�����:��)�T��t���m��dz7J�[W�)��P�ANT���S�Ԉ��_Q�*�0��\^����_��!��tŤ��Mq1=�\Ov��?o
��K��`�����:��-�F]=Iً�/��f$�_���h	��5�$PT�-+P㳻�u�����&�{��B�� zU��aH�&]E���:q�$����A�������B����<��u�@��g74��6��D�S���7b��2٘�rh��fj����4�*��A�k��)5uݫ�9�M�G������W�@ӈ�&��j��X$}򑎴���w�.�����Ǟټ5Y6�7s�@�ͨ�#F�����y_(o"��ı���!	jb��D�	��#���K���s2WQ���A�ki��3�O(��u�dL�&��͔�l:s��7�:?����}8�����Iƥ�e�n���G��$�xw���D����f �V�d�/n�I�1<5���2�]�Ȋ��1��~'�C�M]�a<�5��J){`{Ph�f8����^��\�0?�� y1��� tYrVЮo� ���[�ἰ��x����ּ��h���]��%�m�>�)��T{`i}�2��(������A������N���0F�j��)k�T�>�~a4W ��_�>d9�T!Wv?X��>h�l[��*����`�-���("*w��w��D���$y�h:7#�ʏ8;/6m���/\9�d���E����fƋu����^���n�I[ܳc�e�cĀ���V�m�Z�Rqmf=��x��<����b@�������p�2��<�����.�J�Sq����p%�lV���h��r8Q&?`h� �����c �_	��鮊���}>�v�Ϫ�'���<rt��j����C��S�!Q����s($�$���C�x����N�1��N��2PY���f2Nk��0^��eo/EcTʸ-��Y�2'���F\��
u��Xq�]���&���x���#!�N �����8�_��x=*	/i��� D�$����+�"�~�r�WJ�s��i|��tJzY��r������Ä���ǟ�~�_�d1xo�d���
]�1�f1C�Y�����p �y؇���iAC���$	���� x������a�［J��Nm�*S!��2˨BUg~U�E��<�!���k�i�{�%8Gn�E	1ߝ�$F�)��)}Ϋ���]�,���M�0��d�g�A)���:�
�m���<:�JM���e�Y]���[��>,��8FWSq)�z����5Y*�n��iMͅC�N�������g�	 �W�F j�ʆ����^�E�[�c8QZe��~<U�W0����m,���8�<rw���e$�Qg�b�O�xX��`�%t�h�����2.~f����Oe��(��О&2,}���M����ɧ� s���m�1���	�*׌��4�f~��aї�����K���pM�͆�\��֬s�g(�@YF���V�;5�\N��{��oú7�<�{�R,c����©[�o|�Q
 l[|������iw\�;rr�>)���>{�@��cb�K�,�W����+IP��C��l���V_Y{���Ч��fh�n�*i7�C�懧]����!q�pp6�#��M٦sm��3P��M+ ��>VV�L�������c�_�s���7��ndV4s��˶[��1��������X��qK�qB��-��,8K�4k��w�a���?k�i�f�bA�X��b�S�h4�A�`�4e�#7*��#>ۈ2���r8\��n�é��&^2�O�}:�mQv_�Lho���V�w�]Q#*M�I��0���jE��� �E��MZ�}h�}�}b'S��}X�H��Г�;���ۣ���'�x�K¬�mU��J��	Ռ&����zz茀���Ýo������e4?d����BF��e��T`����+�<g�V,�kJ�8^��~��P3b�������Z�?|�����=�s�ow��V�`�
�l�Ȕ�1u��.Rb5���G�p�deaE����m��J�	��|�>|�7��Ǥ˧��D�DT����2y�oUd�b2��mD���� )�A���f��3������57,X��X$��2T����4�,ϡNW�raB�Vq�+P��p��a��L��r��P�E�!��z��'�)��є>>2
r�ECV�|o�⹝Q�A�Խ��*��Ͳ�7�z�y�e��σ�K�N�%v�;x������3��xX�?�)��m�Ň��s��+'&e�&R$?�l�̊C��"���=샿����S���MA�o���=dDB��,D�Fc����mE��%�o�*Xg�k���&�3A*|�:��d�З�}f���V��A�x����2{�p-��˩^	k�I�'��HڷG:��B,��	��|Z��{�~����oAzkͬ@��*�tぷ�����I뾭��c���#�?����_��@yM�@����CH9m Fy��C�8З7h\���RJ����,�-S.�-#�~ȗXm2���T�5�8�$�?��Bj{MhXn�B����o�Di��gdb�"ۗhw�+Z��B��ބ-F��]
���B�Vp+�{���s��m��h��tT�WɅ.}D?3#x�&H��Ap��VY�`X��5�R�I�:?�P�L[)o�G�<-����Բ�Y���
�ŝJ����mZ��D;&���m=�`R�:̭�+O�@t�c�7�x���e�<�T0�L[ʑ��q��V��9T�ۣP��E߹A�um��n�8di���ɷ*�&..��`��238�C��>�	�0O�����$�4{q���T0uY]C��-4u8�p��8�Y�I��hG�x��@"]5V�8Q,R�l��N���߳�ۧ�c�ꋖwV�2(lʠ*	���c�+����[A6r�XlP�O�G#n��r_p��脚t�/!���-��R���k��Z�.K ���w����G �@7�A�˔���o�跅�0�%Tl�,*u��o���XZ�������[wN���f.�m#Q��l�D#�����x�J�
J��F(���R�],�3e���+�����5�%������fL�����'��,�Gv����?[}�t�J��W6�� �Y?�,H��yl�8�cY�B�FCX=����h;��:ł+��U����%}!��p g�8��ݽ�^�u��N+V�:��a9�Cm���kD�ZN#�[��w�دB���^���/'��[4ja�YuHd���z0s�L��FS36�U����c����cT7{�M�4?b�m�ۣ�fw�@�?�-���rрoB�(�.��H�g��*����)&2��Oʀ���*�c�b�B鲑<ן-B�VZA�Fv�}��M���k�pA}�OCŹ~/>[�`P������D���т��]i�F��*[��&�l٭I&�0g��m@4��O���������8*��l�~�Qej�A������ُR����������F$ɟȡ�ac��G��pz0t����u�(�y_ؐ��z�J 壻'^��J!���o9�~�Con�������"�������DǢ�53�<CC42j~| ��1B�O|��&��,=�C�oE��W���uW��$S�4O���lzM�ر��L�bkuN��s��\�ݯ�ڣ>Q�=R�B]'n�R�q̨�0^���$�"�֩F�U��p���KU�G���ɵ�ߜ��6yB����Y�P��In��i`K.X�_���آ�x�]*m }���K��������!ڕ�,�cDnfE0��B3M���Ǥzdz[�'�_z'�&�%a�y��A���ǰege��s ��i$��-
m���U�a�q���3�߶g�J_G s��QY'1���t�r�\_a��:���fY��r�"���o�aN(�]%���擳WD���B����YD%�z�Oc�a+������:vl�������rK�Omj�c�U�͕P�ٗ6;�7ut��,S|e���C+�*:4O��#�S��.���+�~R �PG#q��r��$��;e3+-ԝ�iyYEֶ'�k�ix�(��Y�kiBVm�A� @�R&L��oQ�ǿ1�n/��rHD�׽69�?}v�6�Ș/ �
Z���_�eT���}�-�k���W��څ�w���Q�C
<,WҖ�z��r��� �X����a��D^�ɽyh��s;&���
��� Ԣ�~�GG�±oW�̛ _-�����v`\�ئ��B$�v#��%����8�b���x�[�V&}��1�Ԉ���ߛ����#��{?�묂M�X�	�M%¯��+�9�u$V���� 7r�=q�A�p*E�e�]���41�������A�䜓�,y�(h�.ʛ�XiA8c�
 خ�5e��΋S;��#k�2��Zַ�1�T���6	II�}[���7����O����]	�N�>��⭼��~��vc���=��n�p�ٶ��]j������.�d��r���������nll
'y���I�a�9��b�<����[�|u���֥h_�.o�x(��p�b�����c���&�W��Eܐ�y����o�f���!mu��j�VH��fN��.��b!�^߳�K\q�ŪZj_�&L�A�v�E���.<�#H���m)��j혛�EgOx�c�)���6�p?�Hs�> 6<ǁ��a������(�v>�/s( ��o6��qN����+|�u�c�U��������W%D3�����7�dW�*	�l��C/������'�/�od����AS=�������a�����rt��fҪF��sb{���=l�=WIQ�t����i�Lwɀ��~��n|�
�I'�'z	�%X�Mz���,��"ΠKB=Fo�l�l��m��pV�'[f���"�^%�BW|-�Ema�*h��M�y(I��<D���|Z���fj;0؞�B���썢��&ģ�Zʹ���jrxt�^�	J�~5Y�;��4WQS����,�������������Í�%�mI�����߫7s��x����)5��<�-�͕�^�5~����d���N�_un�ع�,���~FP"WH��������i���������O�AQu��8,�~Ky��(��1��W�3��Z��r���9��[ڞc����>��>}����0(�y>����!�:����ɪt!蒈�e�-�t�� ���>|��a~ �Z,4N���7h�687���5������kJ��f�\;��'����⌾��O:k�͕/�vZI��(Gh��m
�%�5�f���@�Տ[J�l_�����j��H�n;�25aݣ1�Ӗ[19H��~n��� ]��gЎ���T]��I%~����Re{�q~.�;�1H�c�wa����������?�č��Se�9]vS<%����u�N�VO�84��P=��j�m�Vl� ��@��}&� �Nr>is/.�1|�� ��JomҰ�Mt7ɧz����
H�w7}���`��<]J�;�ש�2#�~�$Z�������PΛ�Gd�#��O�dS�6p*����}J�77�ҶIR�[-H�@���ڢ�#}u�㎛�m�&�`�(��9���o�#�%���C��J?���j�c~��d��v3�e��Jĭ�k&�PIR�O�M$�Y8�Y!��j;���1i���?3�$6Y�e0�B���<�����_��^g��Gí�^�2��h�5F�V �ׂ����44t)b��;S�=��V~%;��fBR-#�`���/ ��*����	A�6c�Q	+a�isOb�Of�&P�&��hu�q/1TP�8=m�J7���8ƨ&�m�b�P��)́(��� ���PK�L�Tcy�I���x�ѩ�l�v� �	O���}�޺��{M-�q�2%1c�^��h����:&����o�41�(|5RY����g�8��i')`��eU`�q��<�����h���Ŝ�$��>��,F,���j�P`:�X鑊���:�'��d�j���̮����9��D�P5eʎ�����q"���1,XY;�L<j�[3$�Qں�^�	�7�0E�"��a��a���Rln��*�ۋ���F�����(��ex�5w�%��x����T}����1j%L�� ���R�A���������M���LgE��h�ِ�n2��E��뎨�d���W 0}�ȉ�Y���
OvX:���MJ�^�Y��9����T/s���Ә�B�A�(�Hj����@����5T@IOEŧZ�{^>���6	m,�Y
��s�n�X��4�hz`8�V���5����7&F䪧Y�5�RP�$∱�@����'����(�;��-��i�&e���}7C;�$��낂(�C=|S���QzyX:��Q����|1��J�//Ǿ�\���x����"�1^!Ϙ���8rN%{�L�g�@8i�ƈa<���e�Џ�O[�Ջ��9h���3D��O����0FhXo3on|��j���-������R��u +z�1���_Hۑ��Kն������@�2�WGq���T�)�%�����jG���"�+A�������4/�9͂�l�>:�����
�|Y�n˶���r&ґ���>�H:��Au)5-Zy�$V���4S"�{��6Ktm��K=���?��B�@�k^K���G0�!1h�	a��r"�<�4a�x����yŘ?9yH%�t��	纶x�Gi��,Mg�S��u���3s��h�]A锵~������N���"fc�@�.�U�?�\�TU9m�ȤysA@�"��*^��/�-=�m&v�	s�g�cQPܙ��f��
W�
���k��p�%���X�`�a�p;w�Z��L�p�B�ҽD<�`f��S��'��"��b���.�T 3�i|�3֎�)ݛ�ׅ�A4��"�T�6X��żpR�Dw�K��Ć��t�1u@%`�c�QB$%����]�fut��	M��ٙ��]%E����M@W&��;]�Zl's8���/��.����\%�0�:<�u�µT������S:ԡ���i�JMY��:鹱���6��Sh��y �T5���<W��� ��`��_�\L�.R	�j��}2@�gz)[{�%��]�AY?S2ʧ.˥�;��V������;KTp.���]2@N�%6��*��N�g�XՊ	e�m�j�n�L
�e�}�I��-S1MD������V�(x9e��W����r��ﳈ׻�Px�b��'h]�Ȣh^�]���o����댻<n�&,0l !��p��i��K�R�Xk�(�~��$�Q�n�'�h�������i�}6W���@_���R���p"7hp�%� Ur�o��̐s�_�����0�����/e�P��%wFbft��zK�L�y���],�Q��!۾�7���u�-��>3��B[�D%�^"������0Q������O