
module fifo_decimation (
	clk_clk,
	fifo_0_clk_out_clk,
	fifo_0_in_writedata,
	fifo_0_in_write,
	fifo_0_in_waitrequest,
	fifo_0_out_readdata,
	fifo_0_out_read,
	fifo_0_out_waitrequest,
	fifo_decimation_reset_out_reset_n,
	reset_reset_n);	

	input		clk_clk;
	input		fifo_0_clk_out_clk;
	input	[31:0]	fifo_0_in_writedata;
	input		fifo_0_in_write;
	output		fifo_0_in_waitrequest;
	output	[31:0]	fifo_0_out_readdata;
	input		fifo_0_out_read;
	output		fifo_0_out_waitrequest;
	input		fifo_decimation_reset_out_reset_n;
	input		reset_reset_n;
endmodule
