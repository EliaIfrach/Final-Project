��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S�q����]�jJ��:�YpbpfvE���������` !����1�W[C��-;w��X{��Qg��Y�;Vp�߾2��š п��::&]��Cm�[�)(:��f�ޖz�i�	�AbN�M�{�r@9����ūHa�|�6=�۠(Zވ<�T0��*�?K�^ψ��ʹ�&*��o��[K�β�T�>��� �� �\O��G���̚�4c��!�D�*gcH��L�J�v��P)�� $_}�z�BO����5���4�R����4^kQ�G��m����!#�"�)���A�>i���1�2Sn�-��#ۅ,���j�d)�&~*�Y! ���$�##/֫�F���^!(B�|l[����I��@��CՎ*�����C�`#��$E�Tv#Ot)=-澾`�_z�T�qP��aP�s����ZHd�h��I�s�C�[]I�U��(F�&�p9�+ֿ·1�4h^�$lL_p���+�l���rm��<Uj?�<�ʿ�Q����b���+�+,��c!f͎
&rp��i�o� ;�>y����7�b�A��t�xL��=�Ɣ�C�"��#��M�-ɠc�\\jL���/�^�5��2N�!�&��Ǒ�t할��_`�U옲I�.,�r��QY�*�+���e�����~��l���Ɛh���8�	��%مE�r>�K٣���zwL��:.rQ��o'|�?�m�IS�5��	|X�mX�6�؇3BX*��h�p8�S*p<6�D���aZ�	�}.��{��L��b�+�k�eBJ�Xh����5'��hF�r�s�w���ٽ^$e�\y��P��Hcb��_&Ӫj��jxi^��M/&C��E��	G���-Rhi��ؓ�1V���U#Q�$#˞�}"tn�;f%���Y)����^��f3��N	�$�Q����(b��b8�=��?���Eb�,�>��po�G�V��r\ߣ6�WD6�_ߤ>)ƣ���Co���d8�|�U���s�׼ޭ�yWG�K����7�ԵVQIʶ��N�����y@-�b:Z���î����_�3�<��>�;�d,y�')c������~!�7\�X6��>@v����$�>����l��|�N֧d��F�#�'bd��5Z��?2�:��G+������BF�|��%����O�v�j89A���˵du#{Yb�C[��? �*�����o`�7x�ޚ����O4�ʇP�!)�@�I��SVS�B�|���� N{�+
D����$�ǬcPg}���|�f�l�L�������ʪ�ē�� ��vr���H'6g�?�ٙ��:?,��+�V� �k�&��A˓8����?�����z�����Ȗ_$V�؃��A����ٌu�^��H��
ǰ����5L���ؒ�3
��k���
]|�(���E3#+ �Җ7~�f��hє�j��4������lJ�tJ#\�b}e@{����X��������G#L �&w������𶔢�*`ԣN�ޜ"�J�#dS����̰L)A=ڏ�Pl=�ĺB���k�PT�6��c/g3������y�m��S�Xdd���2�����~�-�9���L-�O��c	)�`��8���/�>����e}���WLA���.r�  b�b�S��|�e7z�:-k�>P��{�q%?�Gje;������d꺁�%"O"��_�
$U�Wi��ꎂ�n��.Iv:�G��>f�o�b=c�����8���fsůZ���0M��]^�NB���'@��	0�|n-�5����:�})v@�7T�ah1A��$�����p>�S�z]R�������57	�2ͬ�/�q&<��ͫ�yDR� ��~��$Ǘ7Ӵ��tD�"�;����c����zD��@��.-�����2���A�k5iƭ�J�>�M�9�rv �ƽs�A�C�5L��m�Su0A�ckMDKL�b2tȯ���ّ�9��%�_v�
���@1J�at_��mW�@���%������s���U��GfE��u��6gWɁܻ3h��F�Nی!��=�ލ�|�q���e���*z��T̋�Y�;�<��#��d�j�k��)$Q(�ݠ�"�-��5n�G*ۏ$7��NX�O����{���{߅���q���+�Ndm�V	�.�-u���w�lh�?�c�+��hڳ�i�ݒL����
�����\KM�KȀ5?:�]r<��l!�$K�f���7ׇ�s��/�p��%�ʧYS#nd5G]\�� gf
N��iD;k2�.��N��$���G�J�Z}&獵o��8�D:�;{ȌT�r�L�X��ϭbw�u�Y�Aq����ߊ2�;�Iw�Y<1 �+�m3T P�%�����Փ����(��h�"�và�B:=��~��֭��p��#P���؆{y�8���U����b�mAW>��]`�#SbjGΣS�0�X�Z�e�EF	x)S@�7Ɩb� ���C��m�]'ϻN[��-O�Q���b�"<���QL>$5���f8�D���D��>���Z�A�!w���؅P� ��N'��Fz�=�,e��������+}$IL\P�R�lm}T���O��4�O(?R�}0[p)�p;t���C��Te��;bP�m��y�+P���K;��kȨ�˙��g
}�<�R1\�)��Is�ީ��!:ﱒ�eKu9V[�rߑ�lc��ݛ