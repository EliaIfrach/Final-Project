��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S�q����]�jJ��:�YpbpfvE���K�b�1�n������<��-���H���W:��O�#�1&�:��>IyЁ�7K���/�t-j�Zkf���d՛=��r�IC�\�x��,��8u��/i��,K��"/��.�4.%9��MC�t׋%;��=��oƟqXM��}t����F�y�w�9�������r�����>ŋ��ًk��~sNwI�n	���}����l�?#�����@}}ԭR�cI��匰�""|T,ӴrRӬX���Qf�χ$z�l���c��?�y�G���υ9b1{w� ���&G�o\I�98��'N��X�r�*������y �v�mr2��2��.Yj\n�(�,g	a������
�8� ��������d��M�q��<+ C��B98�0<���8)�a�0� C\��SO� �J����V�[���*̲�-�s���Jڟ}/E�)��<KΑa(��~M]uUJ�ZN����a�n��~X��������D/T���X5�a�D�S�SY�I�ְ%%�<OM_�_��e@�[���p�^vI_���-��%*jO������
��I�l�\d��}�eH�������7dM�6=j됧0>1�5�Ε���A��"�Y0c*O?}C/-t�����Ƥ�j����ȋ��\QhwO�P	!�#i<��EN@9��Eǅ�XLĐ�y��o>
�oDKd~
РS�,�-�U��V�46���;3MI~ud�a=,�0�����a|�\�`	<�s����ˁ�J��$>��/Ś��	l��:
�e�Wz:K@Sj��՞�&=�+�zA�����H=Ի;��X��{������HѦ����4��I7n���
ȫ3��6B;�xA�^���~�c�u��������f�(V�3zf�zԉx��ܫs8�?u �I"���*�*������nq�����;1����;�>ښ*��6F 1��P Z���H;�#���{������~��\���(����k�E�Z�����L��!3!dP!
c�;"�2М�߼���ז��c~�*2�⁻<Epc�%���*�}۠X	уeɣ`�+�v�@L�����p��=.�����N����/�����Fx8��-�5;��B��+����vK��L�'�Ay܋�y�p@��x��ڸ��
�WY[]GF����&S�s30k���Zl�s5�*K��H�Ƚ{ʒL�}����Cp���j��c.�J�ĩ� � ��VHUFL�`�mX]�/Z'L7��Z�f��<���E�=5Lu²��^��_~!8��]@�-�a����i��z�aם,�Oj6�rR�]O{U5;Kh�����K���vX�'�����#���͉��>6����H}9��ȅʐ;ПGTXh�!&C+Sc���ϩ�'J�1�#n]�iPX��*���b�j�'euv�$��sQl���G'�-2���*�p��zM^sk(�dwS��"���Y;7�o�0��R	���䨽d%~�༓�Oٷ5���}�EJ �&�$����o�����x%���n�<�(�\xz�,e�w�c�pe���_҆����3�D��c
_	����'��8|O`��_f��y����4�@�C��+����>P��y?xC��wR:qH�jW�J��gO���!z�x�:W�K������fR�y���V���f�\�S+� �[�EC-�����[�_�c4l8�H�V��K���?r;N8	�+|m�eG�P�L$�k�)A"Yx��k�����F����]��Z�AkM@rG>QM���	)����mL��#�?�@����B@@�+�͜��J�Bn��q>��5w���!e�� ۙj�'!�ٓ��k���C;��Y� 3?#�~��b4�0O`�I�-��F�$�����)j�%$.��_��w\鵵��:#���7���Q��&Zp��NH�MT]vq�)��-�H�p�2_������C 5��z�P�i��t��z�����ڿ��i�a�����;�s6�噾k�6�*n�l����t%�!j	l����@-)N�Ӯfx���<���E �����y��̭Ŕ���%�T>¦�)��Z�m��m��k�@���?��\/_]��9