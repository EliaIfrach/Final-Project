��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��-�ro��i�����/�$��ci��y�'f9*�����(�"�5��>�H_��T��B𾥘����DН�E�H_ϧ��o���s�-0�p����^	�'{K@&3�_^��(̕�e�_�_�p}7ewFb$�����Cs�:�<��q��ፒV�y,7�d�,͍_�X���͏�"��U��5��sd��J��a�����M�`��5S�Ғ]�@�k�<Tn�N-+�<�ZNP��p2�aS%*A�oXGm�Q�+e�6N|ə�#�E����H;�w6�B��s��>�6.ջ
��7���,p�ؑ��@������Yt1�7�<e^�h�b���8{���u��Qf���`gbU�[�=-�{fkX��/��U�3����Y^>CC��)!aF�t��Y��b�MI-Û��1���+��K9';"s*��q�Y��@q-���*ͅ��J����8/��8W+=�,�J1����g��-�3*��:��J1�Oۺ��R>���F)�L���M��,�Zvqqke��-���cWφ��9{r���h>.�l�p�b?����f��)��a��ɑ3B���N����2�L���Q���s�f�8у�ճ�q,DֈE��*��ъ�����ԐP��yA֕�?g���ղp��!G�P�`H��)g@�L�K��Ź 8������ɻ��631��K�\�I�/8Y��D����Zr���9|>��"Z���o[|���Ibk�����>�h�ۚ)�fhb� �P���G+��ωc���r@��N�O���@̎�vJ�Y%�����Ҥ��Q�~3ɖV_�/D���qVCz*
��4�KfI��V9�#h�J�d|�tZ��L����س럤��~���������E� ֊R���8�ؽ��-�Y=�G�s� �vF1h�A?MG���`��_Z9� ���Wʈ���o�j�YϚ�̆�l��ǹ�Lү�_�@w�Q�B������|��X�1��eG�LS^�"�"!��K���䋃4m@~�jN���&�\��@�;��Y�K1��={_&ۍҞ�<)�	���V� R`�������L�g`�c��@᠌n1�/�����r�����>5U�U޽��\Fa�`�����`}�Q4@Ff�9UF�V��l�%�,�b��&t��43T(��q.~T�s����Ţw���;࢜7"`�!�z�Z�m�c�A�&�D!�T���Yb���AM�~����$��3#��z��K׶&zڅF�����)�G�V,_��Ǥ�h
m����p>�)�cGI�x{��bʒ��u�uY<)�|��ݑ.�ҿ��W��r���}?X�BL����;�
fRT�g �FRs���Pՠx���!��\k	��d��$�J��1T�t��z��A\i��Xz
3/tS<���v��u�T�e�(�?T�@5�\x"+ޤ��(���w(`��2{wpI�^�X�Z��R6S� QU#9�sUܩ���@��]>���I����e�S�r�7�5�F'<�&0P�ix'/�f��^ncYeJ���(_[A8�r��P:���o���^$���������J���P�3�q����r�T�$��[����q�5
�4%������q�`�W�/����ȯ����)�6�V/�{���p�c��_�{�� 6֑�:R�sC���,��+����4I��o;�8�q��D��W��0�w>C��x�K_.&�o�����Lo�K�%1��հ m/��o�Ś��~*��4�g�B�����&w�,Be\Ъ��/�S
���gd�|ku@/�Q��[��
�B���0���"��>U��]	��m(���z��cH~D�&~A�������WPZ�")�e�G�a��M��%�_g�x]`� F��A��4�F8�
��J�&�wSڃų�{=,�g�����U��Y�*�)lX���������l�v���/��r�X~i����7��O���o��~uCՙ?��0��PA����o�_��W~�"�,+eT#V�����W��<�`�3��5A�X����qy��pҎ�����9'
#��j��֔޲"��� �����a�&'�K�����jT����EO~E�߁�ISmA�g�oud��Qٺ�1~wv�"�E���2)'�)�;G�Z	�����!c�n+q�����d"��6`�2��9�y�=���|�@���!���臼�w4��jd*�m�r���� ����JOYe��]�������jFW;���p�dk�M�q������y��
��6���F�pc7[�{�M���x��hT\�� Ow=�3��@?څ���-���:KPr�8Y��}m���5�(�od�����Q{E��Ϲ�`��f�RqC�+�%��dbfDmތ\��i@�x�-K7Ც�Hr�B\��>���@�[�ձ"t�7�*������w��f�ٚ%��$���pm����v������g��ƱExZUw��W(w؟S��rۂ}{�+z���8d��p-�!�2p,'1�+�<|+��]JO�9u���G6�I���$(pE^�6��K;������)�Uݡ���w�W���Լ?�W{�^r�D��c+��/Qm��@�����>�����+�4���^�ˀ�I8��>�SZM��`�݀�G�e �6!m�����`��'���ckNw?�:�M"�.L+� ^�(�> ����E�6:��ӽ����Q����yV�juB'����<��&�8W�A�몍�����;��H2����䟉I�P������L��������[���A�����q�%d��>�w�_���4�Q��o發�4Rx�!��F�ƕ�Purȭ�c��1w��lE&,��%��L;����涂�F�=�}�r�܅JU֖R���-��������C��d�9�r'�(����������^q�G�݈D�4\��iNY�����r��7꽵uXas�h|��$�R��?�#t�1�	�
����K#���Tۙ�V�����!�.A_,�%���m奬���o�ŋ��u�D��o�`��˓r�_�+ӹ49�`We�i��\�&��
�!�W&�6���
/y�sG��H�_����ޙ^�w�;�i�E�6_?�͂�YU�)O�����!�S,׌�)UI�u�/Mu����i���w+�$Z7�qz�����H�l2M�O��a����I ��f���$A��~ҙ!�Qī��}&s�2�@̓J��̓���'c	ҧ��\u
�ӳ@<��+�[avb��l���z��G�X|Ytv*'�Ξ2�w	nEۃ��IL��Fu|h|"���3��U	�V~����ݒKW��&0���Un��z�������)=/�����3�#�1��wUA�����F>_/x���~Q��FyD�9�62�����������:�����lAp�D3��UQ�9��`$��d���o��PV�a��^�g��3S�_ �+.�B;j�q��)��`�q�	ȫaw�7�&3�2ɖoewV���#�lBV�����o&�fqO�gB�]��S�ϱ?C���[pRk#@��(Jݣ���J�_i��������w���p�Jw~J#��ψ:��X��&M�E�rLi��6�����7u~#zJħ��i����8[WD�����o�H��Jq&���8�B�O�wŕ˖�����WcC����j>N��{�.^���@?qr�wl�g���<̕�y�	�D�l*�f$Hτ�=Y=v��+�ۡ����(��_T`v��{�I�{��/���p ���� F�9�+��]I�{A^��B7vd�1���b$;��[�k!i��|B�Ɓ|-��fn&���A���� �\�:�s�R��g'E���t�?���%����P��=��?y>����NN8���uֹ$5��OI���5��/1E�	A�m܄�~1�B�!BAsJ��gQe`�Y6$����p�Oyp�!h��
O��0�W�`�J�R Qn�.!��u��?����t��-��$4rO�|�C��sWft�J�N���%�6�fX��M���Q����@XPSL��(���nd�p���&q���C)ӎ�CB! Ŵ�N�,QXy��s�u[H��u���w{w����d�r��Z���RM�pP~�ԃ���Հ�\�1���������R�6 ��?`��P�-�4��1㧒j7�m|\������T��"$N����h�0]F�y�$T�}s�X_QT���&`���X�/I�/j���j��,!�qLj���grq��ur�F�WV�"Eƕ��wu����dߔ�/���H�>N��DU3�Ƹ���t�WPi ��G~�}_�]�'�?�sT��X�i@n[m�)���]�7�=*� �M\ǫ�l&-��B�ʛ���yw�tdͱS�
�\�Z�]4�M���	��(H7Y�9��]$؜�`��Α���uْ�������<�`���������q+@B�I�{:�q`�s�����:U"*7���<����v�+7V����6k��*(S�`�` h����m\#0 H`��͈�D�ۀô�}�f���z0��l9o��Ԟx�)���Cu��f�UbI�zVV��-�A�gKt��\.�F�����
�)�+V�o�.d|�����Ɖ]�56�h���
;����:P�\�X�y�7dJ�&yŵ��fg��b(Z���|���j/4��,����/O��.E��*�ʹ�9��1���@"�aX�R�m�!�7�|0*%�a4�. VSP0X��0υ�����J8d}9S��!:6]#W�w?��<���ݞKgk�N��1��D��v��Q�[�g�#�n�z�u�TV��E����x�/��k�/�t��R��'_�����~�	�`g>w���ΛÞx��0;-7��1.�k�~<C��!�y�e��U�QL�n�Cmԅ��}w}�v,���L�Uq�nQ�fS�u��A����A��	#������Y��h�Ո��XL��Y&\P��`����������sL�b*�[9@��'I0��&���e�����<C)��%�����H�?3��x̌�5[V�MȘ`���^9Q� >�:���:E �A����٫H.�۴T-�E&�uCQ����품e>39,��E�#�P�w���Bݺ�p�3mҔ��D���lz���{�o����{��:ܜ�x���D/�����M\4=��˷���s�!&	�Q"�Zr͙�R�XrW\Ϛ���r ��Qhk��vE��&�Gƛ�����?���7��V
�|}�یRr_֎gs���_�)��&�����o[�@!ht������Z���G���L=nE�������,�>HLe[�(��4FϺ�L�$Ie�`'�E�O(�	-�_����ׁmiw��M[0;�1��ܱ�U�r�uiu�s�У�4��/9�mȥ�d�R�Gٟ���C���Nn_c�Ƈ1��K�E��S�ӌ\��i��x~�u��\���>��#��l����J��jc�&.�M̟'�M�����Q�m��&�:��Y5����?�3ۿ�Ǫ8��RJ'�=ł�V"{���JU@��Ʌ"��n��vG��N��9�D\ط�������#��!Pã�vdg"�n$�D6�	 ��!�LM$�2��Y� �i��<�v��q0ܺ�$�sV/6���v��둄ߣf�B����"(ں���¿��a3q��i�M���0�nSr[��".9�+�}�l�\{���כ<n�����D�X{��y�qw{b�����m}���{#~0T�弿ؖ���P��#�irZ���@&.���x��<���(��P?&4���?o0{&Gȶv�'��'e�|�3
6�O#��c$W���v�E/��e�W�sg%h��5`�p{s�`����,�No62�q�Y��]tf���M�.x���B��s�|97������W\�R�e�"�>���@��D<>��[5�R'�P�����#F1�U-����u��l��P
�� �Қ�=�[�t���=[7�r�'�mE������6���aW+������Ľ��`�:-��!2��N�����9�bb��8�h~���ڧ��Έ�A�6A����,��@X�8���Bк'�!�����A�}����9K"Q�E�VQ���o\�A(j����]b&p��+�Ә��޺�D���:Δ���}�쫷9��p�A�
&aO��g�	�=2i`8`є�Tʮt���92%"���o����H�D9 2��%2BT��N���:�VG�wm_�Qy�&��Eȼ����`dz�����|��^O��� wH;����
�
��
H 7�Kw ����Q@)�%��lpT]�4��"�~� s��2�e]\ �<2�r�l�@X����u�4���2ub��()ZZ��5x�M�Pe-�5Gq[�	.�m�YS ������ �G��Iw��� Mu�q��L�w�E�-�;�7�V�U�S��1v��nQ`�x
'w�����aGU��I�HZ�]5�K�,�:�D7�9�tO�u�ȾW�Y�����`~�k	8# ���;ڝv�AY{5^��2*�HiQ��2R�h+X^���Y��\�Q�qE�G�lV���U~�"��>�Ь>�THѡ�u��!5ғ��qC���'�Kobq���%:KNU�����%bW�4䔳�0���KU���k�� kv��?���h���eT�x�^�֎:�����DηX� ���*��{p�9����Ǯ�0� oA�VJM�S�"K�r�]��,�C�]��cEO�:��D;�-)��	��ӧ�e����-z�愐 �v���F��͵+JK�i��k�]��8-�����E�V�n�YX�4����͇��d$�	/��Ū�MK���-��~FeZCOW�"9 Ԣ����r.Xi3�Ͷ���nd\���~�)�����"�NQ�)�I|r
Iw���~�i9���y�������}t5