��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
:����g� j�Qr�")D��m\�5��'k�);#�\(/��!.���D��T��������Jq�c4���
�Pc���$;H�����b>Hh4�AL_��T#�:��|ʣb<�n"��<���f4��X�~�8����fV>��;nؒ�K3Y�G;4T�b�a8C��d���Q���0W�*�;���VU��t'� :�9�u��#@�>�����e����ퟩ^���2���s�N1I!m���ȹ��{J�������p�` k45�?��cp��{jj��7��S�(���>���+��\H��b�or;n�Cz�W���߾,���<�5�j���Z����K�/蓦�O��/�j��]�v�+^�;��n�;��A��=1��ɨ	���Kj�2�=u�I��70�ý8xtQҺ�0H��x����|'�z�l��g�(AԸ��[Sٿ��N#����2z�5Q���ֻ,B41#r�J���@�5��r��O���:+ߣM����}Z��[�;��}�YӉ�A}k1�-1d���Z{v�e�ଵ8d���T�W0�O����3�~�x�ꎼ<���<�\���v��hs �^�{o�qWˉK���x(�Cd�,��N�V�b��w2����Ez����F=��>F�Ck����qMXb|:tvo
�,�Y>�`b�{0�V>OƦOy���U~Y�����h
.��ȿ����ˤ�Qؕ	�(���l`�q��L�F_��T��*���hm:,lƅ�ɟ5���du�P��W|�X}I��P#f$W��≼�yM$\Rp�6��%��I��'��I�H�'Zǭ)��ݿ�/�G.~�����PEzG9j���柍5���b�C�s�NH�?U��t�.ly����;�I��ݧ,�`���~s0��3m4�{'lrW.0�օ#���JZՌ�F���"�Z� i� x��\�����I���C� ����jGY����:��vm�t�J��>��pC�"����1w�+ׂ�	iD�~:�k�qO�yg@��o��^8#��߭M�IaH��#Tk�D����ȑ*#Q��Փry^��_-�`�E��
�ͽM���YGܙ���M$��$x�u�ix��
T�|x�_>�y�9��Q�ֽ�՚����Ӌe�l�PM�A�]eb&:��ֹk�R�������ޤ1ւ����j�G1��Va�%kۮ#rk�}�$�l��E��|���|ʵ��?�bM.j1��6�������=>�1}�_���VXo�C�$�\�|j[�p��^8�]�5���6�v��N��L�d�}5?8rrYi\F��6.���������c��V�<uTV���O��x��I?G��_D�v?�r�"i�=��%�~v��Q��d�I<<R^���;�č�]U�����?>�tm����Q��<������k� ��FUn��.�ķv��X@<�(�������b���{�Y����WCIQ�4 A��w��/����V�B���&\G򰡰E�T��'*��љmU6Z���i�B�e�i��~O��r�5k�!�sw���f��]������D��lj+X��qK��q�S��}�vؔ�ɶo������!}$SU0����M׺>xo+�m�X�j@yX�\}������r���9���͌�.���zn�o\��rl1�Ms��R��d�ɣ֬7`Ö��H���l�_�s���u����cj����βi��ҵ�^���td}���ڕT�vj�ݝ�%��x�;\q�x��:3��±�(�����ղc�k�))���>]#���B�۠�(��b�A�p��ao�39�)D
�R ����+a9x*��t���I�_�C����&���[�ξ�k�9$�G�4�~1�F�;�o�����a>|�"LY!�a�'�1Du(�((q�G"�f����1�
�?�#b�����&Ux���k#ӽ	+��yFxo���T��p��v�ʸ�**��j�6���Mq�':���-Gx��D���j���c��;t?w�$-��M�e˨ ^$~���σ��`Qt�gLZd�v�j#��-�.�U��;��SϽ������6��:����O`�8MK�&I~�٣��c�ҵ�� � ��;{=�@cJ����w�$-y�Q|�#�|𓀀�
{AJVU�;JXl�d�=�p�3U����W��BD���[�Ъ)�)7�� ��Q���{{�ۧ�p�
����bh�B��b�
���YԫW�=�U���e�~8�Z9b�zT���=u�߾��j-�97�!���T�Gߕ]n��l�ơ��T}\�#�.���PAj�kX�<k� TWǄ`�N;�	�]"�*F��\�h�HRȽ(N�@��"�����1�v�Aq��'��#\����m��\l��v,�Ҫ��Q�1����`�4�Pj�(��U�A�%��v�/����Z,�y ��b��B	������n��f�P���|�7����q��Ԇ��@}1���<������^�������%O��GS��:�,E��1�Op���$v���˼c�PPT�R���'�o9b�7+�5��}6*�1�r��,��Av˃q[��8�&��|�XKRT�B�]եJbG^�3!��Nh�;9"��FQ\�!���絹4��L��@�l���L����j�w�þ��e
3�pSM
���A�
���@�㕂�{�e���F�3��|2�ޔ�/����v���8����ni��Mm����@�W5�R�A�X/AX�bdm�h'�)�=!�`�Xu؋{|ׄn̜� ڑa?^a�����ȝ�2R���ч�GW�
d��C��6�8���4�,�Z�:�!���J	3*�����|�T�~�?��:a`~G".u����y ��V�1t��Z�\N�{Q�~��T��H�}���ph�D3�m`����u��1��Ӽ�T�$]���5@�;	U֪��c����خ�8�wȻ��b����>Y���z|�G5���̭�.O�F���wE��3Ͼ��Z����RN�#�2�x{�I\�s �Ow=��;w�@�Zy"+�>Lx��XPn=��@��G#N�&m�6vFG���M]��דi5�"��֞��/a��#e�$�uG�k����c��*ǘ���3rKO��y�i3�%vL@Y!E(�Z�z3�g��_jFi ��eB���(��	+�?=����/�*Ou�z7�	`�$����������v����E�R~��/��IQ7 �g�^��|,�Z�W���.��T����9���u���Ь��l�}(|��/%P]W���MAH���E���؀�g��vq5��hN<��)�J��R�c�_#tN�!�յ'��`���V�X����f�t����3U`���V��a�Fɟ�0z��!KgO����N��݄�Z/�]l��?#���6��9�wա��T��g`u忶إ�I���~�J XR��w�r�[۴��?��%�<
ny�Z���͕-r�-{��M��?�r�]#kzRT�F'C�&�U�("؋�=�Gϗ�=_�R��}%{ۍ+fx@�JjJ#.(�u�!�����]�{�{Z�sMQY�(7_]�����h��W�JP�FW���ՀA�.�K,v��k�T��^,V�1Z�X�P���ͅ��C���	N�4Y<db���939"L�\z�~��*U���a�vuX���.�^�˙�!�O�Ծ0*�ec��I���H���7���~(	��J���1/v�]��KB�)�7��������@g��Z���B[B�b��� ������-�Guě4ѧ���Ao��	?�<��~�
�Y���q24�e@�7;k$��b��BB����:�n@L�«ª7���=�K�y���>�Q`���1]�ƅ\��E]9K\9ǂ��$$Aަv���ci[9�p4���<#.��J��0�:�ü��y8yK[�2�qO�Up!!���~1������[�q��p���#�_ț��O�ru�mH���Z�+����i��T��o:����-mߴ^�#��n�� %:�f���c[���!�Yc�m�Q)t�o�1>�D�:$@�e���/���1�C���sP�6�x�����V`s�^ݓ��j���`���e�O��:�&�k[��աzb�������޸��Ŷϱs<�}�Ziu#AG�2���Йs��D�{�F�<�5/Tn�����6i�R���r�X�7(�'��D$;>���5��H�#c��g��W��ϚF�a����[���D�\^�=����`]�ƚ���m�7pU�}�67ɭ�K �E��~�e"$[ã;'��Cr�����V��s���k!�3�j�*�[����)��5���D:�A�23����n���eT���;�/�\'�8�*�_��0��/����N_�W��9�8�F˼�ꖯ��4?$��kc؏����2�?V$	��^Ux!>�B糶�,G��� �##�ؽ�H���P���&Rg�e�O��=ibh3g��L��aїC�:F%�'b��#G;���@!q����8��0e�V����6��ބ4Bx�(��+R�� /T�|�.VP��U���	�9K#`񓙔�%VVE)&{.W	3�H��������2����xجceg35�+g^g�	�v���?��n�O
u�4S�s=�Z���]��!��0�����W�9A'{�>�v	Բ����5���{2�Կ�X��1���K��gu���0A��.R�9i����� �,+�0+�8�\_�>6(�����V�k�I�ё��U�e�Ulv
7k#eO.�R��f��*���nq׋�r�k/�]�yUX�O���n�]�}[br�/U�ėX���uT�d^e�5��1��!8��`D&A�����h@�u�%Qå���Ԙ� g��y<�1ؐ�c�J�������-�].��^�MB�\���ʵs��%FY��)�V^ �Jg���z�7x	��!֍�g�;���3D#�=����w�\�FP�r������@��3~1@���hY�%�e0ۢaq��h���Eng{�_ �jJ):IC��Y(R�v;��q�~�G�w6ꖇEČE�HVg��9����U련Օm�L��$}h%!TW���@<����`��X� �$Wq҂�b��{1��6l�!=r
B-p�1�N��'���٬T�L[�VDQzs����~����g�q�1AF0�`S�=�Q&EF,��� -��&���j��O��_������NSLOLD�4�Xy���M[h5�P����k�
�������v�A��=ж�;}Γ��׻uF��Ε�&�O,���*���_��{`y铹�3��y˯���k�
~y5}�U�<]|��E�������c��Ġsѧ�K%���d��p�uh���G�?���������T�ģ2����I ����X�����3�iQ\��ݶҗ�f��~��U�����z�W��H�:�w�+}1�rP'����sQY3�1���7p����dO��uFS+�W7�� ��$�[�u��y�����MO���\r�!(L,�F�uI���-e��j�=��!K]�K����8��j�9�VI�u|Iq�\� �JsR�E��f0Rڽg�kl�1Y8Ũԗ�ig���"��ᤤ:�4a��+��;��>�1.[=��Zm��m3������y���I���u�R6�NS��Ɨ�����(^68�kO%2��"�j���G#*6	����@�e�/=�o��3�����n�*N{h6�� �Oٳ���)S��5	����ĸ�]#}�$m���J���U��W&�b�)H���+��Iu��߁���R�=�����c ��U(i~��/��ܴ*5��o5)W�D��#�&��>�2�U5V��O7��I�{�],�17�%���	���1p���X��,�~�@���CW|� kNF�N���`���J� �F�E�Cne����H�C������wJz$�A���P�0�p<�!����
,]c���3��Syf(�'E��� p��d��.�P�-&�e/�J�W�SUV�x�����E�W{N����������[����-$��@�'y?P��1	�tD������F��E�S0���f���<:�߁��G�F�G��X�7Y�ǃ�vx�5�L����S�\
�큎��7���d@37�eZ�"��k��i��/:�[Ai�P��z����Ր��>���e=�� �k��\a�����eC�a#%�"����︳\�/Bud�5�z1Ķ]�ةU�Ht�M��rs=����<��
��Cg��W�_�����q���`����7��M� �����fo>�|ZB�)lS6<��&Q�����UvZ�������j�#N7��R؟2;2��C>��N���/��ך;��q�A{h��.���q79z�8���/Ck���B|�`n�O����H�8��#��Ni��Ͷ����~m!b;�e'&0*��/!!jG̖&�,9���JB��Nre�R�GW��%�_��uУ� �n7"�fo.=6���͵� ��ƙ���ſP�8A�c�_�o����W�Uz�o��7�SJT����������ő��se���Q�������%-l�z�Jc���~_�u�@����|
��Zhrb�Y{��
5ێ��V�Da`���=c���״����u�6m�6,^b0n�)��訷�}t��P>��ooCe��$�0;RPt���T�^�@`\�Eٸ� ؅{eT?�Hܰc-�g @ Z>��<���~GDM��[��FhS9����5��(:�!�ߊ�+���������?jM��WXF%n~ߖ��NԒ?)2n�˿ԡ�@�}�v�(r�wEP����V������w2Bqq-�e��-G@�f��� ��1�.�j�wX@N��K\�V#7N⌓0��ou����Ӹ��C�\2��G밹����w6Tsڑ�0��(Ii&�ϓ�&sö8������I�6چw$v�Ԉ��]���26|�ͷp �o�V�i��T3��yq)K8�'c�PL���b�=q^+�v�eil ���#��}�&�+ř���e����F�ؔ���*lB6� Z(跈f��Ho�
65hE���IM;wG6��'N�H}G!9uM��4B�_H��0��;�
{t��=QG���y�V�����W�D�d��T�"[�[j�>������nk��,��:���M�G	�=0�nj�Qp!.�j���m-���Z)$�m�V;v�t�n �%ȷ-��I�4j�i��:�!�,�"����>��t�p��d7.v�K�3�W�4�׬29�
�fT��޷°������E^��p@[E]T���vWsƘ(K��YC�-"%���#�� s8C��xT�z���#pO���*��jT������U��`������/�����+�
����؋_Ck�9�.���Q�<�"��/�65T^�b�C�UV&2jJ�aӵ��_���V��呇E�c��`΃!=�AKz*D�\ai�ZJʁ���K�
�>�/��'o����S���E��֓�A\W�E�F�F�b��ު7��c(@���|�UZ���p��kJE�0�'�}��q"+�*�-�Z̭��jog��ǧ�x�bC��v��5AJ����4��!��,܈<�����(CÐ������� ��Bզ���)�wV�I��2������O��d�m�08kv�^�X�x�2-����'&�	*��K�'x���s�E�d��8�"����g"?����j��
���v,
�nk�>koJ���h��=Ƽ3~:i�G�{/�U�V,u����T�8 p�4�{��A�փ�����V����aE}w|���SY��TR��x�}%S��q4#�A���l0%�$�����D�g���qSF��q�3��vz��Rz(���m *>�����	6o�H||��{~�����(��'L;�L��1���0ɑސ�͍Б�v�N��+�,����YJ:����y�\�l4)��g�wm^��y��`�%�f�AQ��.��b��\��cH�i�t}���Q��D�v2�@��|�)e44�V?�V�XvC�^P�h��@u��ǂ��#�U6�дUb8��h�il�t��m���~��J�ZB�j�)��$�X��}����G]/&FTd��5��=H�Jv�m���m���mBrW�ݪ�@�?��M�/EF�}0��}�Gu� ouAD� #2-u����<Oر��V�j42]��v�K��N�9���I��ѧP��a)��l��3��;*�Z�Ս��qR�gD�`EW���L�)6��L��n����Av�${V�	�a��{ϾJ%�\���UU/��v�U��='E�n߽�ү�P�%�rb�=��Ѹ�)����� ���VD��ul�|��1���0+��8�2����0���m�����B�d�Ҵ���	�zv���7��^�;�9�n#��� ��']L��~�96�n`�=Q��jG�L ���%�1�'��g�b72��'�?PS�:T����~d#Cs�zPI�3Rj�j����bݥ�g!���И
���y��d�imz�)��d�&���P��52�#�T�|GT}+F��U�]Ȕ�,�d]��d��0 ]���L#���r�sԸ���@�}^��I"�]e���Gɝ���z�P�2d;V�§���߮��0q�ޚ���HVyPĉ�mY��C��k���Pf5��Ȓ3��S�¶���F���o��p��F�yA'��U��V#�!#���/B�|��#z�Y�;�$��"׉X"מO<�K����3���<���F�6a���5���Kr�(�ڪ9���7e$��A�Q�\�z��"�Wc�Al�K۩Ϩ<_�M6۰�Ft�2" �JP�� �"^@�!��)�S���BT��㡮�����L�.�o�KO��0�j_����n!H�as�K�-ғ޺~�p�!LG�]�)y������v�����q�>V\�v'M$� ��E-@�]Z������&�o�}��=\��EDq���H�E������I`�S0T�"���@|RQt�)[�DBH\!ղ	:��Ϳ~�Z`��}TCf����8��q�����uُ��Y_�f���a�*��f�l�G`��3���K�Lʟ� �m����!'%��ӛ�o��h�2���?�O�0��!��˘C����U�&n�V���Ƕi�d��*��������a���M�2�����ޭֳr��7yK�bM�l��R���?����'t�y�<?������FV�4񞔼��eѣ��b��g��dq��A+�gJW�#lH/1[�B�\�.��bs[��v]x�?}6�cxa��l��zl����1F뿊�֨9^E�>�(:!V2<nf��yPM�c��(�!G̚����y�q�Ư+����:~�l�TB���f!������Ҽ��-� �qt��}4/F@�<+t5�Ⱥ��2���� <����ȿ�~27#�P��㩝�1[%��E�֠����P?�;��tc�Y���$/[�Nc�]�8��d�y��|��̝�@/�Z��w�S�ˮ>sn%���7y�h�~fgB��w�V!C�we&��|�#~�P�t~≻��)�X�	�8fIt���4��H�p��!S�VN�('}ԙ 7��e!]�"� 4ptz�j��q�g�eb�FR���h�K��l��w]�6�<�Q3
!yIK>��������V��t!�ԣF!��0s|���:r�V"J��)W&VVAr@��"�p�]޴� Ih�#X8^�р��3��r
(��;6��_$�'��F��(�:�^���(��4n��R��pwUu2�·kD�G�;�-+ˡZ�>�*�ck�nZyY�K�MLkx���c�2���|�d�'�m��lvT��&D��ƒ�T�mO��BZ�����
�ďd�R�A���lq.eq=�,�z<	��N�_W�� -��iw:}���Qh$;���D7���k�R�ol�ū �\���ry���f�&�(��z
����<f�ځ?k+�ˈ!��£�٨�k�dŦ��9ع��9�JTl���J���{o��϶��|�x���<��F�D�_ۯd78$Xg�T]���M�C�}�����3{/�l�V�kz+��"w�$ٳ�ۉ:�]ST�\ߔiGJcT�y���Q�tn���
"3W�����UK+*w�]��f-"4�c��"$����F���{��d��i�I&�n��3ּ~M(�T�UϦ1L�a�W#��$Ŏ���7:ՠJ" J���IgA^�sڀ�jc��^�c]��"F?�t{63�R!'�2��,�)���/������( �]'0/�}eF'3H�<]��Oގ�@a}���C�͔ۡ��v	Tz���',��E