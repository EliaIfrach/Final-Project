��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
ܓ:�6���О�d	֡I���������]W~4��vqVzr�@8&$���0��;�����+��$6�0ma�·�j	���1��;�?���I����	�$�Y**���~T�6�bnH�l8���q^%��Y�ܧ��.g&����K�K"F0TԔ:2:m�ɺ���ʓkR���~]/���V{q�$8z�9y�ZTV���saF�͗�CP>wi������[�qГē�IZ($�����{�9��(�8���c �$L�<#.�i�/�=�9]�I���f�F��k4�`��%�$Ixn�%=�Q�;�z�*�qA%���|�%I�T.V�6~U�T�:��'�,ا:M��pM�ܫ>uɛ���B��sG]t�!l8�V���K���~��Jf8���Vي���d����Geܟ��a<�C>
�'�$Z48�����`H���ح�K�����
�c1�1�U�1I���A$�9�3|q:lZ�k��6�Ӥ�Z)�d'g���As��T�-/o*G�c��p���*�]��e2�{��-yD*���h��0m�B+�K`��#Ϻ �<�*�D��ZS�����pcғR��������6�� k\�������uD`"�����u>M��1ң[�;	��Q ��*Z�l�K4 $Ȱ���������"�mj�?����q�V���0��r�Z�7�p���7x����� 7sб(]��5�#x�<���Vo8�j6�y�+��>�N؇H�+�5t��^�(S���!�����z0�-ch"quY��������h�]^P"0_���a��^&q�4�W�)��L����O�:�[�-�#;���#��L���.TG�����m�!� ��͘�ǀ�8�0e�w5��I��n��a��>V�B�pۆ�M&�����9��UC��#>u�*�����W��01���T�|L�$C�]G"uS{c�hJ��ϖ='贑������T5�]~��G鑌��i��7�E��0ZT���v��=�6�JƯ�*��w&Q��.�Ljhk��\U��w-G��=�����t����;y�Q>�T�!�b|�G	"˛*.P|���ܯ��ߢ\&����|���q[���۹�W6bBK!@(�؊�X.�3�Xp���p�ܐ�w|�P����J<�Rtl+�%M:�1n#T�F��z�/C7 /\�z����F����}���$�YT�~gN2Sc|	˯W%�Zr������Jg�Y(Ć!��̐SU��v�ԭ�{�^&A�V�o���A��귊����AHqc�W� ��鶙�����F��̿2&���E��~T��f;Q��^���ЗQAtNoȔ�!�d`���L���q<��ж!1;6��LΗ|h���_3�L<�li]~f<�zy�A�Z<��>�2�&jɯ��%�a窲]�ɪȩk�5RVH�o��{����&�{��sf��r��nPm�Y�5Q(R��W.�J�nV3l��64����w�V95L��ytڟW��쁑�T��:��Ԁ��]*|�w��Sn�����˔����x�|qH=�y��|��~L�c�܈��&�_C��lg$X9ނ2c��asb��ړ,6�%����B�paq���T���������]Ƈ�DB2�b�	O��ߙ��s��m��B�T�waZ/��6WiT��?H�~��>$�Y⧕|��G��/Vz^f��r�5���ۆ�HK�x��Z1�ݧ`K�RR��m)�+YķB,l�Z�˸�67d�,�f%���;u�\��5�\����d�R�%��Gl���g~�$F8z�fk�c2��W�-vj�/�Vi�Hum�*��W<-�;WRt e�GZ����8�N��?�dE�d(��d=[D��M
����mQܹ�������D�є� 	w��_J|�`��Q���3��f��䨶���Q�T�U����;x2 �����GF��n/���ǟ���+SCS�1T�++��{�q��38�5�'ZR
@Ȧ ��*�H}��g��Qp�4fxwpPh\�x�ij@x)h*
�v�hc=��>�� Y����4Z��6�kN�f6/@�t�Oyy���)+�"�eeݥ�k�
�Ym�4���qk��F���X��[Iu��P�������z�_`G���?J�i�6�!��`	�j9k�C�5�ѫ�������|x!%� t��Ot<������]�G�Q� �Md���X�HIwh�r�|9 8�
� ���	CN�^�Z7w�e�A�������ߘo5譫�F�܋��\4�"�ՠ=���D%O�ٳR��� �o"����Z���*9OFl� )+9�My Q�׹8$�g�oX��2Y��]���r�k����hڋ�i�/����v���!��rH X���+�z���t4�M_�M�N�g��C�5�ta���q�)���b8F)J�wEw4g��^z�xs3lݕ倵9@�ɦ��L	��	Z��a0�"��m|l�����<Owt�6o�F�3�ו,<£|��B��;M���C��a�ur�"M�Y�������ͅ{��^m�ɖ]gW^��ja���F;f掃7/�匂Q��@IW�92wd���	X���2��s|>kL;��:���ݒ���P{FFV�ɣ�*I������$G�R:�.�u�iΦ��^�b]FpS�e��<�j����J���+0�ȓ ��(Y��)I��(K�}尪�P+�_��tO\� ]�������x?�R�%�e�UL��R0ڸw�ꙓ5�1!��ԛY�DŒ[`�s�v��uC|�2�?�Pү�p��!��=�4��*�\j����e�eyI�8��� k= �xI�e��������wg��<K��_�ߑ��׃�*�~�i�s����J��pE�����&�;i���:��������[��)�#�s�g���`JѸu�_���R��S�N^I�fhca�0m�V��-����/]�ӟ�8w�zCiٮF���t�D��Ua��:���8�t�'��|,�ܖA7�-��)!��^��Y���=ʡ��oh�|���Ջ5:�7�,b�T�� ��U��i9O�/t���q�n���e��ċ� ��'�J�碄�M��Z!���
�E�:�s��~����P�-�d$S���go�[�vB{6|jQ������>����z�5��NY"t���n㳆��`��Y�B�tM��3�v��!�U�V�0���f�K�Rx�A�8��߉���Q,�tV����]EH�ؖ-���O�/�D�	�4PH9.�"P�R�Ձ9 �;����:: ai��B�I�H'Bk�,�!��;��[x�-٬�#��T+;�o:&�Hĸ!`{����h�v�Vi���tG�%��5�ͥe�de�.�|HK��$y�IȓR%����%_���bq���_��K�����Cݤ]�p�#�� �[g����'���ǘ%��7�q�����$�֘ڹ�/:�"<�n�j� MO��i⟇�V��H��Y��ԷR���S�.�a�B�>%��b�(�P�F,ٔ�S�+S+gY��)y	��eC �Q�DnC ��tQ0�ɬ�\ٺ&�o{�1нL�O��{(f�����ͧ�C[#�od&�~,���^�C׿�-�7�`8��i ��o�����*ҢQ�+�Fr�{|���:y�fCݴ����;��I��F� 
�F����s���2�,�@�PO���,�A�Q4�A�*C�OĆ,�+t��Ӷ͋�ႏ�Q�Hl�s����U�t�<nz$�Of��\f��W��ӯ!�\[�ɉ�ߎ������f�QJ�*��B��	���o��
w,%������|j�x�����0��L���S "T�h՜ �̑M�d�Y?i�� �,����s�>6T��ؚ@>�ڿ�b���__T�B��'y�Z���L  B%x/-A�G�R��ٌّ2}m�
�|�Is/<��2/�bf���d?�IW��6j�m�E\RL��X��z[�h������Bu��X�X�~�M����l���e�8:���5��4�͡R1�����ؖ�.�u��������,�[(�v��Z)8��k�H_^@�@��� ��k�-5���VB�:��+.�8z$˪��2���r���7#��$��k��g^f�>��s�yU���#!���\}l�J�]�^/��H���J�hrӴO��i��,��޵P�(�t��a�=��Bv�9��c�f]��g�E����C�d��͕#��Q�%p(�����d�F�l,��8/=|Y��{T~�������2{
�c�����B���v̨s�L�\���\��d��`��$�Si��ۉ��bR�}���A�TΚW��Yq�&�"���xv�j�*@��`A�r�R�Ϟ`����/_U������#���0�/9'+T�8�ep�bӬ_L�ğ���(���]yU�t@���p������\�軃�F�1�W"P�u��R�x�����U?�U�f�`�Mx�6"Jt�	B��+�e�cvh�+tt��˶����ǉb���*(��\�>��x-=J�� (�	�[5+���O1������ա�a��g���w�G8�A�ю�,�Lq���.S�Ќp��B���ay��7�\gڰ��bwk.�#+k?�x&~M.h�%g�N�2:�'V`si�	 qQt� ���/4}
�<�b�2�L�N�����������ǌ�3y�MMsT�Vf����i�es�NO �����j9#;j���6Q���Ƙ��X�����J�h�Tf���(�Ф�tc��	�/��E��Ν�1 �a��uJ,W���^i�̭Q�E/VG�� "6M/��Y!���eWh�\jJ��xt�9+�/��W쵲�(���Y�<�eҗ
Z���d��A9*̝5�|Ǫ� �g���#;8����������f�b�Hoc��� ��t#�nH+�#V��b3ƾ��C
Kf;��5�g��ء(c��猯�8}��d�M�Gk�ڂ�l[��f܌< /�
�1h�¡�A@�yRh���|?%򻔸�m�>*�ʃ5�Y#%gK��Vt+O�|fm�6�n(����\�ƚ�0j9aF�-#�����0����Z!�P�b*�&��:�׾�ֽ�m�����L%���W�L��S�
�.M?�1U���鬓�	�S_й	����7��q�B�i��|2v��t햄8O�_���c0���M̸n�����$[�D�.E��5'�ٌ�:, ʛ�yOKS�W~b4N�χe
�����,ޫ��^� B��p��q@��G���vWD�E����*0�"dæ�M�P`���e���r���TG�,ʲ��E��Ic�JK��\����T�� z��fNW�zM� E�Q{8'�c\u�}�gA+��}܆�o <U|�O�5����-���W�jX"j��<��S6�6 �֢�$9���}�#y~q��s`� �ն$M���A���\Lt ��;����XcٙͣK�C#����8��nB��wV��Ǥvv���F^qס��7T��FfKc�](�QH��F z=)��L[�^����DV�)���T"��L�7�ծ�n楽����)VCz�k��qC>u{m�o����E>)�9kw������c������-E=�f���y9>�6��e"[ Fb�t�bܢ*���v�{\S���ƌ���*F�}��7{9RRj%ΒHăM��D��M {�L��\�9rL�L�5��ziH�Su�d�"���
|M�|�N�g&�0UX��eϯ!��0�d�~.{3Iq�-^�����({�cBPk��gm����V��g=(-E�a��s��wz�}C醜z�اAȈ�w��Nh�{I�KS�����zU���;�㼊s�9����N�lzŜ?����6d���M%���֢<���{e�����ȩ?�%�>rB��H�
�D}~bK���?�>z���>�v�<�6}��cf��
ߏ\#��!x�W�0�.�y��_���WS+�����ġ�V�'�}j-Y7�$��������A�F���[�z�c2Kr���O�y b}p_J�
��k~�]���u��t{ey8����GE����Z�a���j!sxO� ��/��>�M$Z�b���X:l�Ϯ&1ۡ(�G�t�<buO�I�`J`X�����q�N}�d����ߒR¶��'��[!�Sr`��s%�A�y����Ǯa7Rτ%�_b��U�lF��8�PաX?��2DQt�ρW�X�ܟ�:k/��ގ���z�"r���i���b�P�(9�z�ܞ̈́��װ�*I�U��W&3s�y	i�0�,�l�	�L����J��V[i��i��ӣܡ��6�rŸ��s�
n���� .$Am�u�7�e\�I@p'>y=u�C�~]~���vK���9/�.�<���,"�֞�>8ǽ{2ΊWw�ߕۘm��9���R��w��!:nɟ��0C����BΧvF��,lH����%����==n��%e�W�ْϢ,AZBֹ�X���?���F�;FƤpi�uZ3�i��'Zf�J�-("�"�����Kt�����(A�����#O&�O��#Mߤ�����s�L�E<�71y�δ�c�?�E i��v�)�z�E�10_^�������|6!���j�3�s.�)tSDXq���>�ii_VfBʙ����ތ��m��ֵ�׋ѿ�6!焪ara͏0ɒ�g�Qx��؛]9���<vV[��?� ����k��R�����R-7w��\�����;y*��[�l�[��!�[%�A���W�=�`jr�S��V�����F�G�<���}�W��Z����^��.�еWi�O'�8"�Y�4�SKqyz�`��?P��	D��r��eB�$=��"�$"[�8i�EZl�zs#�W��1%��6���=����p�cW����j���� �t�N͈b�⊅,�5�` �w�!�<��&�3��j����6��G!��lc���sF����̵��5�8���d� �K2�u�?�.-���%���b +��Q�:���T�-���#�w�?bՄHx1jV��n鎴�&�z�X�`L&U���
����_}�s!�3�F�T���\�ڈ���S� �;�md(��ik���VE{w
Yt��(��I�*���7�؉���#:�:eT�N�@�����SW),��W��}��v��ɱ1�W>c{1��#ݔ2�N���C���[��������~�9,˿Ko-���T�?�z&_r�����O�����f�Z���Tq6t17L�.�TI{�'��M�dH���p � @�B�!Se,��:��a��X�p�&�����+��A��G�a�\l��P���5cLF�&5D`f5�ܚh���7��N'��w˛ �rq5ɪ|f�P���f����247���)��A:ru�V�A�����q�����Ve]�i��UM�������.$ oQ�xtϗ]��L(�_mKvK�qkQ����3/�9i�1S�q����^K������3�P�$�.�t���|���%��uN_���3	��k��'��s�zݼ��8A] ^��.��p� )~���紌9'�����v4��n���GШ�X����e�>Kc6�ܨM�����*��� �!rf��ݭze�����pft�.����sFqj�k��U��0I��
�|�H ���k�%r_Ķ��#l���Sz���	dC��:�E�HH���a[fv?^�@q\��K���"�47�c�Z9��{�ޛ�A����e ^�
�|�5зx���ޚ���^}�o8� v�����n�z^�s�x���%�^�)�����:OTɿ:��b5qS<	�D�>�����n+�
/��X�|���]��ܭ��������]D��� ����[��T�<��ю>*��s�<�l:�^B�c0����<� �H�NF�S& $��A9�N��&�������e�p�.��R�� ۃrvwY)��:`�tyoi�e�I�P�0�%T3C̈A�8(l`2KÎ��1���1My�F�P��#�B������+
:T��"}ꎓ�I�c�&k��P�u0��w\�L%��֋���|V��ëd��<<+���ep�Ij�A{��c0:$��ᾃ��l�����z���d���n�k���ԩ,6Ђi�A������sዐ��+k��ʌ���-���x�����=1 �2���J�������$U�G���E�D�Q�%��}�?���}�_s���Kl���ƞ{̈xF�Ԭ��x|�5����v�lg\>���d�\l��޾��0L}�)QA7�s�^�/X/ap�P ��ӊ^6���w��Թ�{�;M.
�[0����7Z�TZ]ASl�-��H���0F�qR���N3$�ʟq�a�/���h��f.3�PAwm�Ku��
X������u6�x 0�BL;����`�R%�³h'ѣ���K!���b���!Y��f@t����q�g���ijD��$ [���qb�LFQ��j�;���� OXj�{�t]G��Æ͠�Rcv��k*���p�ҳ���S;��?�w[NZ������{K��IS'Z�٫ ���7^�R�E��4&���c��W�"�B~���}��0y�KX� G��/�+�b�](A�~Y��腽���-�K��;�}��,Op!^�4:�Wu$�R�7�%�,���|o�0`��C]GC0��Yx�7�(���Ó޲S�}���=��҆�����.�����V����-��9�������]�TJ�,�I��uH�3j
��9L������5�9������żD�5ỷ����Ό릏d����|~���Um,�(�M���7	S��/��� e�{��'5A����n<�P�3�z���	��
Z(��HK��C<"d��a�Y�֩iG���f�D���
�����v��+؜�%�e��ǐ	�^F�s�3��'�����-%٫�f�딓 /ם^�d	��'8�7C ,��͔���w�%�d�����&���(�˟�:�8ݤ�1�`�8U N��+!�K5÷�|(a��k�N�ݗ���r��Ibf1mk�<�������Ͳh܇Gl:ׯ�*�%�P�����$J�IR�eJ���#���W��g�\��m���#�oJ�=ǒ�t\�=�XX[��퀴X�U�C�b0RqcX/#f��2��rkTj/�7b>�4)�y�PF34�Vw$��G�Y����W�[��rL=��aK��;3ٰh���,�1�и<�a$r���|['�{���yȄ� _��S�Ee��-7�'\o���9�{�o�$�r������+X�0��Pĭ�G��it�P��r�x^����ߴ�E���M���|��"D�xz`�OS0K?�2?)Z*J/��ӥ��Ө��F&�"�l��c5"�� ����:�6�����2PGK���`_��<��Wb�'�]���k��(B<1�V�=m&nX��p&!�2�EQ�l�뷐F��H-|�lx���=;K���n����J�����T�9���N%j���7�"ھ��lI�БA=9�}R%VcX
�*{:��Glu���g�T����%.�=!��~����4�X��'bck]����BBx�8�L��G:��5>e�KMB��tw�P����zq�<6��^B��әe��=;�4��Ֆ��q:}���D����G��sU��)E����[��hl"ǳv�6�d�S���:���f�� ��_�p��i�q�d�z��)�PePk�sī��fq�If�:Tta&�.�6�P�ԝoa��)�G�P�Q̀W�b2�77���]������ڧ�Ko �9d��)����� ���у"���Q7���p�����(�8�?��)� ��ܒ)K�۝��ߍY�����w���S<Č$)��� �E5(+n� ٛ�5�]����L�vgϥ�r>'�W�WR���b!����t�`��>-�nB����tz �:����F�J��DKm4�,��:&%(�j!˄K:�ĵ?����8�]`dk	�v~�ac(sUn~Вc�V�G���R��7����c�nL0<���R��㷕����a�z0���A��#�u�τ��X'�V̚��=s�'͛Ҝ�U��(a�HK.�w�t#.�y����2��C�gnS�����h�v��n�lwz�h��z;]O�^hʩ���(�s{^g׈[�md�n�a� ��@s{��c�F5�.�&%��U�8h	p��ŷ����+����ϝ��?d�����9�dl.��0:�3�`5^�InZ)rwbĩ$�%xB���l̰wQ,b�&�(���o'^T��L��BY���doȺ��0�R�O	3y�avc���4=��j8��lֶ���/?� ��(��h�C6�u�HD�L8����
�x��e�G��ـ�T�$Shmn��H0$&�[��ӭ���ֶDU�!�S�O����	a�,�j{:��yӟ�ˊ#f�h��	����1�?��k���Z��f�n���Rs��"��93}�_��Ӂ5����:��َ���{����{N�O���<}y�W�W�8���Jf�yR��N�uh��Zx�8i�W�խy6�l~:"��F����w�U�Æ�b�|��xUuJ3���[Q馊v�
����Jd��b����#c�S� �P��6�&nsV��ؤ!�-�YN3r��4��>K��O�,�������
�?�M�[�~��f��"��*�)`��`}����z�!)�jZk���^QP��b��JY����X�G����?��/���������s
��)�m$O��M�P6U���8���5 �张:Ӧ�ɻo�9���eͿY�>[	09��c\��@