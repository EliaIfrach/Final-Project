
module PLL (
	clk_clk,
	fifo_clk_pll_0_outclk1_clk,
	reset_reset_n,
	system_clk_pll_0_outclk0_clk);	

	input		clk_clk;
	output		fifo_clk_pll_0_outclk1_clk;
	input		reset_reset_n;
	output		system_clk_pll_0_outclk0_clk;
endmodule
