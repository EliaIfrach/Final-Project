-- FFT.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FFT is
	port (
		clk_clk                       : in  std_logic                     := '0';             --             clk.clk
		fft_comp_sink_valid           : in  std_logic                     := '0';             --   fft_comp_sink.valid
		fft_comp_sink_ready           : out std_logic;                                        --                .ready
		fft_comp_sink_error           : in  std_logic_vector(1 downto 0)  := (others => '0'); --                .error
		fft_comp_sink_startofpacket   : in  std_logic                     := '0';             --                .startofpacket
		fft_comp_sink_endofpacket     : in  std_logic                     := '0';             --                .endofpacket
		fft_comp_sink_data            : in  std_logic_vector(41 downto 0) := (others => '0'); --                .data
		fft_comp_source_valid         : out std_logic;                                        -- fft_comp_source.valid
		fft_comp_source_ready         : in  std_logic                     := '0';             --                .ready
		fft_comp_source_error         : out std_logic_vector(1 downto 0);                     --                .error
		fft_comp_source_startofpacket : out std_logic;                                        --                .startofpacket
		fft_comp_source_endofpacket   : out std_logic;                                        --                .endofpacket
		fft_comp_source_data          : out std_logic_vector(58 downto 0);                    --                .data
		reset_reset_n                 : in  std_logic                     := '0'              --           reset.reset_n
	);
end entity FFT;

architecture rtl of FFT is
	component FFT_FFT_Comp is
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			reset_n      : in  std_logic                     := 'X';             -- reset_n
			sink_valid   : in  std_logic                     := 'X';             -- valid
			sink_ready   : out std_logic;                                        -- ready
			sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			sink_sop     : in  std_logic                     := 'X';             -- startofpacket
			sink_eop     : in  std_logic                     := 'X';             -- endofpacket
			inverse      : in  std_logic                     := 'X';             -- data
			fftpts_in    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- data
			sink_imag    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			sink_real    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			source_valid : out std_logic;                                        -- valid
			source_ready : in  std_logic                     := 'X';             -- ready
			source_error : out std_logic_vector(1 downto 0);                     -- error
			source_sop   : out std_logic;                                        -- startofpacket
			source_eop   : out std_logic;                                        -- endofpacket
			fftpts_out   : out std_logic_vector(8 downto 0);                     -- data
			source_imag  : out std_logic_vector(24 downto 0);                    -- data
			source_real  : out std_logic_vector(24 downto 0)                     -- data
		);
	end component FFT_FFT_Comp;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal rst_controller_reset_out_reset           : std_logic;                     -- rst_controller:reset_out -> rst_controller_reset_out_reset:in
	signal reset_reset_n_ports_inv                  : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv : std_logic;                     -- rst_controller_reset_out_reset:inv -> FFT_Comp:reset_n
	signal fft_comp_source_imag                     : std_logic_vector(24 downto 0); -- port fragment
	signal fft_comp_source_real                     : std_logic_vector(24 downto 0); -- port fragment
	signal fft_comp_fftpts_out                      : std_logic_vector(8 downto 0);  -- port fragment

begin

	fft_comp : component FFT_FFT_Comp
		port map (
			clk                      => clk_clk,                                  --    clk.clk
			reset_n                  => rst_controller_reset_out_reset_ports_inv, --    rst.reset_n
			sink_valid               => fft_comp_sink_valid,                      --   sink.valid
			sink_ready               => fft_comp_sink_ready,                      --       .ready
			sink_error               => fft_comp_sink_error,                      --       .error
			sink_sop                 => fft_comp_sink_startofpacket,              --       .startofpacket
			sink_eop                 => fft_comp_sink_endofpacket,                --       .endofpacket
			sink_real(15 downto 0)   => fft_comp_sink_data(41 downto 26),         --       .data
			sink_imag(15 downto 0)   => fft_comp_sink_data(25 downto 10),         --       .data
			fftpts_in(8 downto 0)    => fft_comp_sink_data(9 downto 1),           --       .data
			inverse                  => fft_comp_sink_data(0),                    --       .data
			source_valid             => fft_comp_source_valid,                    -- source.valid
			source_ready             => fft_comp_source_ready,                    --       .ready
			source_error             => fft_comp_source_error,                    --       .error
			source_sop               => fft_comp_source_startofpacket,            --       .startofpacket
			source_eop               => fft_comp_source_endofpacket,              --       .endofpacket
			source_real(24 downto 0) => fft_comp_source_real(24 downto 0),        --       .data
			source_imag(24 downto 0) => fft_comp_source_imag(24 downto 0),        --       .data
			fftpts_out(8 downto 0)   => fft_comp_fftpts_out(8 downto 0)           --       .data
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	fft_comp_source_data <= FFT_Comp_source_real(24 downto 0) & FFT_Comp_source_imag(24 downto 0) & FFT_Comp_fftpts_out(8 downto 0);

end architecture rtl; -- of FFT
