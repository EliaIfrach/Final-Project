��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��-�ro��i�����/L-�U��lOjj�l]I߫�p3^������_"�'j�ʬn�*W�� �a��;��}���������)t�X�|�r|�~U���;��k��2��%�`�	�c͜��d����/�OB��*$�K�[�>�)v���������~$�sF�]����ZP�6͝*����ĩ�';ɒr����YU�|��#��Yq���65��~�Mduث6z\j���4���E_w3�Cن̷����o�I��Ƃ�G���~T�VO|�θ.YW�9�����I�0�J����r�=fw 	`2K�$]�NF^-F{Ux��L.2OP&~����k2���S�BY�F���iG�H�E��+�%h�<����I�[��G/*/�F��➳��nZ�W����Y�o~r��_�$��\����f�M8D�o�OO���"��D�_U�@��MC�`��.4W��ف�O(��
��,-�h��jn<;���#��'>�鑩�!i����8�1	ZB4J�yY����p>G�����ٯ�`����?C��?��=Y%!��b�IWx+����Q�XjD�I��5��� \�u�u�@n�X�gs"ݚ�i\�X�8�xt���'� �� ��\U,��P>�Q}�������g�]�JJM,��𺪆l�
��z�G�+�QeE"�<���?�PS��"V������FSh�Q��p!�o���M|ln�P2଑��\v����7��e5h����p�C�M"�-�v��4͵ȁF[�=0�$^��ܜ���y��Q$u$���6d�
��"Ｚ#�/��/���34�}��$3#|���2���"�f�4!��Bˢ�mn@��Q!5���SU=��h��qJMr8�q�<l)�Y��Ѐ��������eg�fMV��I-iҷ~$���^e%�����^?⬄�٫%����@(GI��}],#&�M��Q�_�z�-�e�_ ��Ԛ%yQ�?u�S�N:�A���,�Ŕ"	mcߪ�I�t���<�����$"Ϩ� m�/���sZ\�`U���sUF;�Tv�V6wU�zkc� ̡pפ���r$�;�)�%c���) �f�vl�qn�M����jR�g��"?��y�,���D$h�%7k>�AMɜ�ʡ֌/䶼E��G�u�����V��!�`1%�-8X�����tc�xk�"�.�R��ge�|�7�^��w�ă�DE<��P}�z���Y���݇+~����tQ�)�Y9�a��=��һe�g�tV��r���e�҆���YPg]�Vx�45͋m���2�}cϤ��Avq)>Bax��E?��!�Q�g�r��Es��ض~x��b�WaW)�%�Y;��P±��rgEA���F�9�CK�6���6�t9P��!,-��G�P��?��^5��ݒa��٣t6�g��7�w,����wkUTo(�}$H�aj��$��-2���؎4��"��+��%�=$�g;b뙚M�w�����=���Owx6�����b%FA�
�ްT�EͲ��2[Nc4�0N��;�	\�!<�����T"R~ah�{�a]����k�͜7j�Z�CS6S���?UΙ�oz��!k�����<��m���
��X�T�<�|����X����fuW7E�S��&����Ԑ�$��(�80;v��1Ej #�F|�I�ǲd�R���;V����{d��o��lr A� ?�f�ts����=@�P���0J	.��  �i8h�������1p�P�A&`��6��GO�D}����q�!��r�G$���)�Ÿ1{�Z�N��d�t�7��c�=��|��=�R_��'��(���x�G1|<�K�\�=�C��mtG�[8�4�H�m���Rz��W�O���g�d�8����V�{"Y�j�"�>�5�AD�uY ����8��dwZ�]��O�h�{|�%��b9?Mg�Їөn���ZK0�圗N�D�.����D�{��oR�R��F���A��]˧�b*CL�����Y�((Ѷ�5�m�������:YI�(0y��u��Q�����<�0�{������qY}��)\?�i?4����t�}ddj#�+B�W��s�`x�|�e��? QE�.63��Ml]��P@�
G
#ҋ�-�C3ԕؖ�5��VA���v���]{�����yU켴��s��?�1U3��.�0;�`����Үbg��4����=��,��b�s���}�FY>G�jͧX������c�pgD�S� �CXa����J��툪���)��$������t|i� Ka�o9�P}�p�́ڍB�OE�ۂ��>߅��	�����F��!��V�PP�q��G2�W��~�7�M����/�L�6�Cz�vx��[�h��Q��K�|��W�QT�_6���/R�����H�_��z�����曖���tq:�܌ҽ�/k��,v�8�緯�����Վ�R~���O{��4|���yoW����w[q1�T�t: �(��O�༤�:Rڬ���'9�pc*=	Y̸�o����J,�4��"1��p�{u�N�A�o�ƽt��5fH��\��9���(��j/J05Y�;c�Kϟ�:+��fCX�j
��P2���W-L��nCPF_�L'�-������%<���k�i}c��|A<�`LF��1����%(	$����W��,�Qd_,=�X��*B�1�F�͛y"j�"h2�7�p�hO�$)>�uY�@�:˯,<���{Q��^��g���Ȩv�sI��}�{K�Л����CzE.��)�; �ay��sa�z߱��\�P�K�T���t���AqXr���?B�6?	f�<7*����O*yO��B�X��
Ƙ�ُ�(B���W�/��^�<�6U�V���Һ����`bA�Q��t@��i����.9�g��b��]O�W�yj�'���ʘХ���:�Ť�n����a0��'��{-���Ȇ��ٔ�RP^ĹZ��$щ_|nDa���?Y�K=V��r�Ee�:Q��1�b��V��:�������x�sWvKH����E0��5���M�`�h#	T��S�P7'��A"R$���c��om�`�'��LB	�	����[]�ո	��;8�K_����d��O��Mz��
�ÀWf��DI2�
�\m<%����Ê7�bH[��"Y��i��S�"���]A�[� _�\�e�xL���j3��,Ӏ�$�C�|t���
_T�|���4��l����*dn�-]i��ኀRna��R��.DO�d���C�3�`�f9fv@�D!�A�RŸ;(�ƈ����B�.�2���POØHdV�S����9Wi���!����qj,�Q�B�jQ�a��6����^�"_P��������bKH���m�傋°��į.�T�0�x�?l�����{�#�,��lb�<G�w6E
�����6Z��M��C�V.� ږ7`h��`(�5NV���nu���@����u�Az=~�e~������Q�*����}@WDכ���MY����{-Bj��p���ș�HoI��X���(�Zǧ����I�֚=���:�	8�����{�Rw��Մ9�=�NO�D�:���881$7kq��!��Z��Ft�p�V<���Rl?Υ�r����pP������dE����!L��ԧ�j��2/./w$��z� };��7W�2*�����|��2��<���(��I�O�kC��!�\v�zVa��)^H0|�QS�1e&�nO�([�F�}{b�+��L25e1���t�W���mv]qWZy"���?h ��o�`��B�û�x	F ����h��?�1�`߬08�|�Vp���m	 �^�����-��y$�8��")~q(��S��7��>���6����WRf�4 �2�2l�C��&�\1�N~�&gH���F�c�u����p�8�"q��A�����>4��;���ٕ���n�D�Vh�r����kAZZ6����x��5��_˦��I�!2�;)�i��;s����.�a��#�l��S,�_K-B�)�*]����OB�<�u����nv߇�lI�M�jK�I�D����,X��m�3TM2\��u�Y7����N0�������E) �F��5� B�i��s��߂.x�z�|L�j'�E������b���=�h�S@�OP.X���M�f�C4L�L��v�=���/4`�i���?�7J*�{���I	A�� -Wyr��S�_��}�8���M�a膥�"]R�ɞ���O8�X��W�CK�Z�٠�^�͗ߜhm��d��v3�n�����9ƪ�ă�ʶ��&D�yZ_v�A+﹈a(-򒤶�qQ��@�m�FH/�HH)$@!|��b�Ӭ���Y��\15=�而��*�]�M�f����9=u�u�XV�����	j2�b��ᘪߺ�s�U��D����P�L07z5¹��6�K���=|F��!{���WlsQ����e��з��j�7��u/xK��
|_���+�r�͓�a
�;��3 ��V��vZ�,��s�H:ǊE\WI4��	�у|�"��^OF�#8����`� �ɻO�M@4g�4D��s��\4
�>�~ϧ�����o2�x��t�D�'F���'L�&�.·�6���	2d�Y���
>����A(��<l��įT+�j�&�|�
��4ao�[�ȤZ�[*�����'�"��,J�������IM[+�t^2,&�ioP
�X�p9���:���i[d	�-Xu��7i�_Y!�iqE�zu�Y�h74C1���a Ǝ�h3F�#1����R�VD!��x�����ʌ	l�R���hӱ�T<�ԅ���F�&
IѲ���h{[b�p�u������'^}�����#�����)��^c��IYo�=��D,e!����a��׽n�p`S%З��I��\�ۜ?7d�a�/���x�ׇm��-���i�qM�a}`^d��'�p���/X�{�0wqU��!��Q�m�i$��÷;�Ϳ!�4�e��gd�p��֒�x_'5�,��bY4��r��JR�'�/w���`T�_���v��L����^�'m�ȸ�'� F�!�ֹ�E���֟��;f<mi�(���u 9�+�d4*5(4�Z#� ��\�;�g�!v+��>��1�
t��^\�0�ȳ���Q�o��,�Q/�=fu�~!:���lBd-n'�Y������$MS��.�ڲ��G}��Vg�Α�P,<I#��ӏ�����+d���`߉@�s]���J3wuΔm3d�����C��'q�l�ܵ8�D���0��l����׾9I��z����pE�3�v��kk�]5���.b2J�[[� H�{0��X��*��ո��8���%�.ܑ���ts���Z`��|z�B����K�*[���8�L~�VY�&����#F������'�*ْaP{��t��oG^n `Wq�A�i.lW��h�?c<��#�	���q(��
��Щ���Z�(�+}2�Hzϓ;��ӲH�p  ���.�/�"�I�mz=��@�Z���<�̥��j�Ŷ������5b��3��'�HJB�5�2��p=��L>�@�9:����2�x�NK�Bv�l�3HdET��6�Z���M�^�i�f��U�	#՟���0���0�@��2��୛@a���=��2ZߝYXGd ��̍�.܏��6F�B) ��:�����輏����G����Ek��ak�&�������v��;���~�2E��Z=�!i�c#0�맞h�͚�b��2�]������B�hѺ~�Zo��aW+�7�`��X��}*�>��f�Pf�^A��LD��U�/�!����Q6i 
����ݖ6nK q��dm��;�ҝ�{��=�r��ߒY}�ZI�>��zo���sa��!�h�C�-���S�_Q���XU�Qf*��Q�4��0a�}��2��YǸ1\�1"Y'�*��Z1�!v%�rC��pU�)r�Xm�w��m���
�t��	ԝA�yT-��%r�!�r�ʌ �k�
u���_<�t��>U���
鏜sҍ��7o\u���3��[e3�?c'��8{�kH�g�>R���\
��}�Q����;�3L�2���a��o'�3��_/u����rC#ъ���+�I7b�ݗ,G��������ų�Z�� �����f:���x���n38j�VC�޻0�r7��ׂx�d�ƚO5�o���CM|^ UڠP��������jD�J3ф"�Ns̄;9 (��O;��Qb�O�wPb�>;����-?�[
ږ��@��.�/6P��~Y���5�R�xjr���L��O�����Q�����>��-˴y��� m�:���[���_���XC�Y��^�,�r9���\I�#h?�);p���P8t���T����#���
k�6�{�n�.�6  wB��F� G� �BBk��ê��'�d6-`AE���$l�^���ۼb�y#��̿�a��/Ɛ�t���ڮ���!z�/�| ����uԈ[�ˇ1Pg[�C���ZJuv�j��ؚ�6P�CEQ<�w�(��Tv��v:�YA5��z�Zf7A�{������"挚v;ϖ��|Cָ�P3V�_hQN��S*mDI��XD�]6�g��y�+u?�a�o)^.w�p���;'�+�=4i3%�ۦ6@�ᄆ���~qo�-�D���9��za��~�c��z|�0K����oF� �������U�B�Ic
{#j�7�~�o�̲�+�om=�X)�zkm�T��(}7�U��gbcqo��b�է`{7u��z�XR���|��/��l�X�K����2�����X$�S
�E��zs��X���넹�աZAx�����^�{�:s%�-O��ݔ��~�,<Gg��C �G8PW��^��^�mEi��9�G�' ���JtѪ';X����lp�:�x��3���r��9-�=Ư��f�h�� �on�\�=�5�Zj��6hLN�?a��_�r)�ŌV~�Ese