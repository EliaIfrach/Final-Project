��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��-�ro��i�����/L-�U��lOjj�l]I߫�p3^������_"�'j�ʬn�*W�� �a��;��}���������)t�X�|�r|�~U���;��k��2��%�`�	�c͜��d����/�OB��*$�K�[�>�)v���������~$�sF�]����ZP�6͝*����ĩ�';ɒr����YU�|��#��Yq���65��~�Mduث6z\j���4���E_w3�Cن̷����o�I��Ƃ�G���~T�VO|�θ.YW�9�����I�0�J����r�=fw 	`2K�$]�NF^-F{Ux��L.2OP&~����k2���S�BY�F���iG�H�E��+�%h�<����I�[��G/*/�F��➳��nZ�W����Y�o~r��_�$��\����f�M8D�o�OO���"��D�_U�@��MC�`��.4W��ف�O(��
��,-�h��jn<;���#��'>�鑩�!i����8�1	ZB4J�yY����p>G�����ٯ�`����?C��?��=Y%!��b�IWx+����Q�XjD�I��5��� \�u�u�@n�X�gs"ݚ�i\�X�8�xt���'� �� ��\U,��P>�Q}�������g�]�JJM,��𺪆l�
��z�G�+�QeE"�<���?�PS��"V������FSh�Q��p!�o���M|ln�P2଑��\v����7��e5h����p�C�M"�-�v��4͵ȁF[�=0�$^��ܜ���y��Q$u$���6d�
��"Ｚ#�/��/���34�}��$3#|���2���"�f�4!��Bˢ�mn@��Q!5���SU=��h��qJMr8�q�<l)�Y��Ѐ��������eg�fMV��I-iҷ~$���^e%�����^?⬄�٫%����@(GI��}],#&�M��Q�_�z�-�e�_ ��Ԛ%yQĵ@�~�Bk��.���C䙝��Z��,�Y��,_{��/s&�I6R��W�x� �������7�0,m<�/���zQ�2&����J�̗ٛ�Nn�K�xȒ�˜j2������,���l黳�Z����#�;_ c'�Or�i�'��� <B�^#D'����.� .��˨��[�_!5k�=d!��/�	��D��puC��;�Ǥ�*�,1o�s��PK��O^UDO�z� 1Ao�K���㲒D4t�'�89n��Q�o�g�b}?�Y���J�JYXE��'�C���qW��hv���^� Y�d���7-�	)�)��'��ĭ�Pឯ�����v׺�.�%+�YW� �w��1m�&!�JDXK�;����2�D1��W�n(�z0;�ۡ���
�	eE���]�)Ţ!nw��ͲU��^���!X�1� �L�</���-�M�g[��n_7b|a�:���F׃�n��p�{�%�`��I��
�4�P�!�~���E[�*�(��Jqv��#������a�_���=�~3!�c�\�1"-�ȷ�"#��/�<lN��C���/<�,�����{��S�ꔊ�[/�+�jF$*�(�Q/M�r��5����Eйr�:'�k�p�	÷���k�
T��cv�k�j�MKh�˧��k��S�HW�"����u	LP)��6�`��W�F$�L�/���xћ�fc�=�%)�;���*����х*d��/�o���F��.NV@&�8���K����'G`�h.�ߪ��<��S[ٴ��	?�OQB�~�W�mNc�U��������v9�QZ0/}ﱙ��!��ӌZ�Nb�/z�!��*:P� ����;����ҡ:�|D��h8u������R<��T�y�R��;E�͐�ކ'�}��(�h��h]E���p<(�E7��)��z��^�MB���쿜G�?�#�"~ds�Mk5�m��0k���s/�����/
����wT�v�D���;6�M��V��rT�� #��P��L�ߴ�p���`��x��� ky�%Z0���xs��W$)�lN�K�RΡ�Y��?�(�������ĵZ�ڈ9�.݃s	�L���h���� ;�A�V.d��9���6P}���~�j6["R��2���N��y�$�	Vʻd�M��8�9TCUN����O�J[T�|�!�z4��zlI;^h�E��,�6���:\�~+��m)QN-ף���|C����#ń+������g�w�3����b�\T�_�t�*��Ԯ��ů�D�$=�}�Ȉ�V�2�Jy�e�. lVɛ��ӹPA;���>D���́�2��ˌ���~��Dm$�\��� |��%$�����\��PI6��A����i�a]L�D"��PBz���hbb%/	�t�.�����vr�$��C�2,��ؕh\v��n��Es�S�Y����$�&�2�͉��<��D$�[��5�s�L�>�[�!)��׺��J'��T���h�E'd�Ps��QcL���hk�T������/	+��W��M� �]�&d��k��JX�X���0S�d�(���JL��?Z�,��4�iJn@���[o���;W#���bv5�VS۰T��%2!��Z�X$�xi��K���_Z1�Q&���?>��
��-m1����v�_n/�oG��`���E2�!<�_T��р�t4$����©Z���C�	J%��˽U�?��-��'x�$���4�OSO�S>�+��,H�L�ӡ�(l�n���0e�xhx�$��3�IFz��S��ľm�� scq>���o�,:{�	S�Уj���JT]���N풷�}�w�vB1�r+�yP$��\"���B�o鵭�j�1�7�&Fج�"��p�,��8��!���]y<�.4e)�Μ]����4Ȋ��6�B�d2{&�ꝱ���s�����Y�>#	�8�RBd��a�8�D�����L�YJoR�V�KR�NPX�K1���	�Fi����W܋+���g#w�6�<�+��?��M��R'Ѻ���T���ء�>#^�>��UxY���m�u.*K���Y��|�Ë)8Eo��R�RR��M�)���m�6��H��{�f�,�Z����	+ط
���s����+��
�� ��Esq��{�-�Hglx|uB",�����4p��",�,����Q�ox��z�"LΤ�\2�����p{���I,_�fp�¾ubCQ_*��\�O޾ݏ�?���-����78����*��� �-�;�EC����R�u_u) P|����T�;�F�~;�3��i�{��+�Ec��F�Ӯ�:@L���@��k�,�3��b ��Y�h�c���p���NLo+S��q��KO<���|p�s���g��W�4�=N�]/j�c�y����GҠ�6�����Q�Կ�F����o]?�l������̛Xhn�l�\�Y��Luob�:u�r��kIa�֦��Ν���B�փ�"�LG�-�0[�N�N�2 <��}�9�
=�F�x3+�B��p�"��*E�ѩ��7�K�s�|�w�^VG�G��J?¿��Ab�I��,��H	$�,r��
���E�c�]LR��,��.$�my�d�,��W���Y϶0��~���wX�%l<1����W����-]��*�>&bx4�:����̠�W<j��6���n����\+�+c���k�1������H�p.��!Ht j3���n��י�bS�W4߁�C��UT@��/h�+'Z���IE���V��ݥ�% Z��g�;0x�-�b����kyZ-H�8��X�!n���o&O���� p1���B>{t�',�Z�\s��[��U���LN���h��y���.�����	��g���C��a��xH��������FSQ1ܠ���꒎z�l0��%�~r�l�(A Fֳ��dǮ��y��@��s�dj�j3y�̓w�l��|#������Ф��/|��L��=�ѫ=����y���2@�W��N)���mh�b��Q�hm�@A�8:�PsΩ��۠�� 1���Ca�¤�CII����=y�Q�|!?� �/J9M���5�N�L�d���m"5b�D6�lH�V3?�Yd�R�;�CՋ"�^�m#oBx�����-�����O4�����X��%���h�N�T*fU��9����y�g��Ms|�dz៨�)���'T����Y���� �x��w�hb9�hF�z�G9���?Y�ß,�ӻ��2�Vn6k��Tu�G�W b�Z���KL`�p��+� #�M�^t��o۔�/�ΉE��UvL\Vbv��f���@0��@�W�_<���_�ܶn���(� +�z�L��Iv��.iϊ�I�Y���3#�����݄	��LZ����"*o��(����#R�g����z�l7���J�i's�&�T��L���`/�m�v��h����S%�쁣9dɋ�t��;m[�E�㐗'#@`(�+
yp�{t������ �oD����j�ы�䄣�:5�rԙkg9�
�.j�-�����1|[�79���?����xwx�+���&��U� ���ҵ���!��HlK{ �Ǌӝfm��'��Dֱ^Жwh!y�:�!}�z��k�t������:j��^��'�}ȫJ����uJΏ��S���\@a�X���#N2�V�����@bQٜ۫_85M7��I���L��PpI��43���)��x0��b%��+}�[�kg��d@�L��I��i�ǩ��ΓkiJ�|�k�9���yF9
d��
Q�"L@�r�A�.y��;���9� ��-~,1����X��b�=p�@�.K35�z��,�M�h�F,�,c9�-��-䛨�nR^J����%zt˽]�x�w.k��Ü08�ka��C*�k�q:�e��`
T�@�	b;���9������W�Y��w�
�#��4�#����֖���k��ݰ� 㳞����" �0g��l����|<�AQ�j7Lf ����b^�@�������"3Y	��z�hE���A��[ 9�t�FD�|��KZ�2P�h��M<6!�A[oi��Rw�w~U<a��1�hT�J �;�Ӂ���DU*�7�O���&��9�"P���o-�+>q<�a�ci�dwY�j]C���y���:*S��=:U��%u��JW��Ot�Zp�!�|`�k�*�Cml�6��^�������L��^^��vN ���84�Gt�������ʇ�2	>@���~,>�����!8�^2� ��M��!�x�������%K\�5\gP�KL'^�D�_�T���72z�%D��a���h�JN� �����?� ��]�����҄XBq�2T%����]��D(�b�=y��KF�oY�We�<@m�re�a<'"qE�K0���v{�MD��r��	�B�^Y�(ff^��/�k`�ԃ{���m��� ����m�ڞ�9Y�k�L��O���������\ �����f)k������y.����$vc���Y6�2��By^�: ��}6b�y����n�鼞¾z���Y���m[R.�� �]�P�h�a�H����}d�U~�$����m�dR�E-)��Kvw��.T�g�H����{N��4���:��j�;�>N���dt4�mB�$���3�)�\����C�¿;w�!E�|r#kS�A��an0����c�UwxJ�bfRh=���8�0k��+E�f��y�c��^_|]q���!
U-j0{٤j�{+q���l2��x�J�֧�of�FO9�T!���Y����u<3��2W;(� #ӝ"�9�v�'b��d���99aN6J�Kt�eA	?�"��CvѬ2ۉj
z�ݤ���{$��
�*C�>����9��mDlS���s�JVx���0y�K,���0��Kw}'�W��C3���	�G�Cma�"5��Lq`�D� (8,�X�ك=�v^z=Lx�z�0΂��h�CL�'bV��q٣-�§���M��[��fZӈ��+��Z��4lͧ~�õ9cl���L�B�H�{�e�5�]}������H03��_��f�dk�Z^r?8�C��C��)"g&�-Zt�6���$%n��U�uwJJkjP#9fZ�A�l#�4@�����aO��^.C�U�7G&��H��%7cϣ>�i�3K&���m�ݷ��?��
aN�w�� ��.4`�#ު����\�X�'D�Q�]G�h',%�`�ՄP��Am&��@�t
x��q���ߞC�*o��Q
/E(Mru7:��-��ӭ�h(6j��ӵ�W��a`}p�<5(&��R�����WC�������d �HE�zM�_ݞ�+�׿e\~h!x�R�s�x����8R��d�֭��M��l�2k7~ا��ms��ӑg���
bæ�����?�w4�X���Bpݞ6x����,���.�۵�j�@BI��u�����FV[8T;BC��R�Ҁ�EI���- �Hț� 3�a�z`��'�\֎g����mdO��Щ�b.�@��-�l��E#$��5�o�T+�8ga�E<����|r������_Mq��d��+��r&��s�1t ��f�zK�D��������9��ښE�:�Py�Fg.�$Ѿ�9�ꪛ®������ ������HZ�MǾ���
C��$6`����u�`�h�@�h��k[����J:�q}2%����mDC�~Xox�v�6[@�^ {˥`9��yV�p�Ą��RM�
��,�Μ�_��󞓸I���4��K3p�rs��{��c��r�q}l35�=���T#a��;������K�(�tzs�|X�C*	T�������c<_�d��8O���J T�7�_ֱMߐ��g;a+��Jވ�b�� }�\�с��������< 9L�<b����"�N���u\���t}3};�O������b1�V`n3{�d���R���\=;g>[�"i>�|��ԍ(�!�����H�6��)����	)X	t�`�� n��ɀ��_�z���d���o�������tg��Va$y/�d9��Lͧ.�,}İ;7��8�v�V���Ά��eMry!j����eb�%��+1T�0�y�1�?HV#G�"�9N�e��0*����If"Ĩ��"^u/\r�����>_�H�n"�SF���t6c�nn�=p��!zQa/�)�hVN���k�p��D�m�Ժf�6�rݤN� t��]��6�k"yӀ�;� s:��Tz��s��K��7�YϬmyGαg�9�Pr�:M۴�d7����KGx�OٳP����T	S���y7�n�BSkCMAsO0�=9��3�ƭ6�*�����2|x�ŗ{�^9��`����[<���^�r;O}KCWs�U4r��p��,�h���ZC��d��aɹ��y���=�k�{��+��tM�FF ͇��my-�ZIֿx��l:�&S��	��=q���H�92����q5#�M�	���*T븯��K7Ӿ�w��*�;Jbf�>Nl�?�;��u	�[V���5�sqJ��Oh�|~�%�_5bP��.��~�w]�^N>~L�%r��Aku�az���`y�3�S�q�-_5p��p�V('�:��񾧣�U��Z��mV��^b�P`��"{w쾀��n�d�w��ə3�	&�/kt���T��2�Y���Fm����&��7����ڧ�$(�b�#�w�NI|SY��4x�	N�Ğ������Z�bJ ����Bb�ZQd�'�$�T9���W�v���2����7�_�櫬$�Z�7�~���)x�K
Ч�HLs�oB�����~�������?�Ĩ��g8
�nEն�mQ9S%�����RP����˝��iJ�p�N%��4��0����t������)����K�*�؆B `i�n��y�C��",]��G�,��J��;i�s�p^�DՀ�6c���^ �8�����@��=}�$a.�	PK̮a'pA.uwܶO>�Ah�۬*iJSL*�ٳB�����6
a�c�� 9��!.��ֵ_��A�(��j¿��{�3^u�/B�.�}	�]�;~
��3��CId��Z8Nh_�A�U����O[�����������_k�Q�r~�ܠj�b���d�UPߐ���o�.�NS|@�ў��&�|�4<�tiO��F2+rh�u���j!e�뫸#�Ȳ�uW��x�9�ࣹ�Q�-d�6W[T-�o?,�<'��ω5Cz��T�����v�d9�a�Q_<V���ת.t]�^���}�	�@����)Y�߇I���d���0US�p	�y�B��?5�h�v�K�[_
������/�NNŐvE�Q':��ڻ��q�3�5��Iq�?�?ś6Si�KK޽K�_J9Je^��RȨ�� �\�b�z �� Iðs@�A�s�C7� ���X��juw=���U�r%p��� g�-�/�v�M��Q�b3y�����;0#(�[���Ͳlr�?�3�Mru�Zd>zV�=�O��T��fC �\�`���������%�s/ۮC%z��o�u+{h��%�ڰo[��-{H Y]�Sp��EܟηW�&GpxDXt%!�%�[�#�!.r(����s����o��IK\�r�$����VZ; gr#�,H�'e�&�)��F��ʷӀ����5��7JiS�s�9�4��4���A�g)����m�IwO�T�$r�d�,�=�
�c�\U^�}:=��8��|i�ihf��O��UA*�D�M�&gh���e��@�@��N��,Ǎ5��I�"e<��[w�ä��Ֆ�n@k�������pdO;�=�s���O[��±݄�=�qz&��F�{T���x�4ð6���!���XAnF_lK��I��Hn�]%�멓���d�;�����RcY�W���nfօk�V<T������q��C�p,�v��<��gE��T�/L��bS�B�HD'M���%�g�H��K_�*+��0	���Kvs�����bT��7��+�Ȼ��������1��9�}����&�]��̰6���Xr�D�/4X�%�����Oͷ�#�3	�S�/f�V���^%$۾������+3�48�o� �2��V���c����G�����u��@��BogC!�rv�yG?]���*x�B��enOS�tP��Y��
�h;�f�=+�%�����h�
M���Bjb��$ ��w�a#�"�PtQ[��ީvW� �d��1�����M���g��2C�]��u����5�N��:�[do����Q$�k��r��|+��?&.o�
bl��2��Q%��:���d�]�{�효>��*YV���y8dx�G��u ��0�,B��9[�3�tj1�ܵ^�'Y��!�!͵!�u��I��K�x}�����
�w�;�t�s��E�&��'��24LT`�=�fǬ��K�e͒�!��{8�"�`��&�i��o��!k9���Q����T����k�oL�}�G�(�q#:���r�����W����3��]�6h�����T��6#�L��8?��ୣ�,yӋE-J�/�n��e~5�`�g
8�!0Q�u��X�� ��Dt��� �$O������j�?�"��]����%����xS���-6L;��x��@���J�L�?���X;��x�}��'$��W7��ߦpq�������{���Ui�XY��;=D���#��	*�ޏm��x0�+}m���R{v�WA�ZsL))��9N�3n�J�|JGK	M�,�^8���f��{*j�O�Bo�/M7p��ѩk����&^`�\.R�-[ EހYތ+ff7�K~�=t�ؓ�y��_�\���m��5���Q�S��CE"���abN�a����X�O�,�>�@�T}��W5��UX!�jLи��d�������Q�"SG�ٟ� vU��^g�i�;4#���i��1�7!LDn�������&�L�Fʈ�	مb�kOx\��֍0@�gl��=���t������Le%SV5�5Fy*H(��q�]��ejyEo��H�+d�r%O'� �a[6����Tv@����F*��G6݉����m�K�m�y�fɑ~�tm�UX���xa�$T,���Ar�`cr�q?5J�Y�>��RlF�����?�}�#�.� K��g�<��ؤִD:�|���x=�eC8#�.�]>Iah�yFG��؎\H�����|R�U�ܣ\TCWT��BYn%Z��:���0*fc�xE[�"v�l*�%��# �n���n��_�\l���Ze[8�J%�ؒ�u�D��EM���i���%A=�P�ͭ+�x(��Q�`o��2�V�c���J�q ��v�5�� ԅ�����%d�_5.<��Zŋ����ꑜ��p�J�^_��?�Nm5Rpi��.����g{>�zpM�Q��[���g;�$�N��p"SH��n����WSܽ�L8w�t��zdƂ��r	���|���0���X�UE�7�3&/�99�K�Ұq�@�zY�M�
s��i;PN��Mu���'c�^.n��	�E�ϊ_%�B���W��qa��.d�U�&O%�ъ	�$����^���D�1�����kW�H��(�+� �1h����x�ѯ�F,����%�ؔ� @o=*��!kPe�<TU�������p�`���1�~Z��J-�:f�LY���}Nhv���[��4M�i�8;�5�J���S���ї�-b���*��q���v�������SO45��\V��#�K�E������VNQd l�J� �>,[)��a)hWt��N��L���[��r����?��[�ܫ�}��_R3����B%˨=>��H�!��m3�6��\�4�]�h(�J��>�-�q%&2�*����>t�T!?�,%�|N�h]�s�2w�*������}c���T���0���AY L�H.*��oe�r}�c-]sd����AdR_ѓo@�U��l�p��w�u�j���1��p�r���+EV
�i�w�4ז�j�z�0	�)�	]�ݸ��@���ư���ʧ�^�d��w��B�/o� �M����W�c�@�Mt�����;�@�h��ؽ|��N[O�mk����9̎y9'˷x�}{�Gt_�"�w��R�oa[�`���b��$��C����G�����Q��>B蝘��+MN�8��.I�659��yU���'�.�+����Q��:=Ԣ�\�PU$~��8���h�W����i��-?R�u.�YY=��	����0�|i�h�~�����İYoDEU�b�(�'7AA�����S��nv��� `uC����fE\�*7��ۺ%�y�#Sk��=�I�}n�����f�/v&� GI�,(R�K~9�&H��<5�ol���5�L��R�o#�:z��-T��CGM�/��0�n_u �z������k>�Y_�ٛL
����g�\�aj^�לmB�� ���q�mj�
��-�\�c�q3�}���m��ӧ W�jubn�`"�(�j�lEy"[���W�;1�O�D<��{l��Ј;�h�_Nw��蓐H|�?�n,�>RUjۚ���W��j��C��MռQIt8�Qd��p�����equ�����o��ũͯ�Vd|�R�h�_p`�I��V��׆ԫ�
�EHذ"44�*��� nzM���۳�	� x4�>���q�)LC��5@/�O�>�����v��?�S��x�פ���t������y�VkO�U���
�4?H^�f�F1\�=�yb��ll�,ܘj��l�� ����t�:�e�Mm�O9��*���4`
�y�6'&q��{����5�꒪�[� ��|��c���`룩���>����Ǎĕy|�:�`c���Lg��:������L�z>�+��ibz�a�Bmn)+�X�Ù�~�9D��,	���`-���,��x���{�8��&�B�2-�.�Vs웸H+<��?��gF�H^ 7
�$�sT��Z��/�6~�w/�ף���Oa��E
�Z?tN�Ҧ�T�FQ��i�����av�`ɒ�O�{�A���� V�Vj]���a,:���u嵸��h�O�6 ��`J���J쥵Y>�/����������;@���'��*�����U\F��׌�.������������e�7����%�U=��4�0�g�~q-�Txcۙ����N�ѷ����{��^D1���ɹ�n����j�8����ǋ��D��j)�ƈ��M]r���7vxӛj	X�Nd'pk�����~��.�k$7�ӓ�T��F���c�t |�Եp�(9b��}���}�u�oVߣzj�'�ľ��9�x�p�]-F�?G?�������}�N�?������?b�[�{�<!K�Дj�#pG�� C�^7�R�v� ���l0�YZ�'탧�et�!AZ���&�.4���)��I�{�D3ת3Z��N�&��.��lI�s[���T�:�#C�F�(Tz�x�4���`��<�i>	 j����_�ac��/\h0li���OsL��6���ǸS��٦n4Ai�])��`1p��nw�u�ۈjN �s����E#bL/����m�!��R�J[[O����
�b��s�W_�����*����Ìʭb�zW�=|�w�c��}#c�3c�]�����+�Oݪ�C.)�d�p���a�
;"	����Bԡc��
�Sr��J��*�1%Mި(|�}q�e��B�8����W�d�3n+q�\R��z\�Zk5�����q��h�|F=*�6ْ���,�iis`%�p�/J�d��E�Z�3}�+D6'�W&��n���J����TD��.��>Nt�ZHg�]��V�O�tqi�|�ڗ��)dc�0��u���~�lƔ�ɫ���\/�	���X�-b����)�G5x����X5�c@��P=Qo����Z�u;���qa @�MU�.ԝ��� ����,�׮�5t�{�I�-�z��x�0
�F�����!(�I6�����3����c�u�6�a�#e1�$w;�E�r�x�mR�ބ�"�-i��T���7+�&�Ts݀�
R;i:�c��3��e>� ���SA���6�P[�����Nv��Y�� �4*��:�`���1���`-�4�y�Ҷ^ŏ�+��W�z��ϼ���)�Rp���q��[���Q8��_�s7ֹ?#�7��w�׃+"$-�n;+�3��
� ��K+QH�3�Ѣ�i��A��Q%p�\+�����NEĠ�?Wס����0�/�PF�D,?��$M,�e�k�}�Z�GE��2���N�Kؚ����TE�T�\N�2#��{��L(��,G�+�U@Pz5⚁E�ۍ$��x��=1��~�?0�/�FIq3$�����bN��DS�q��κ����A���9ς�'�Mω�M�w��4�;C2=�x�KB.�m^&oo2�P�֘͐��;�30M
t��`�e��w5��<��g��E�8�;B���5e�ñ�'X.�q�DI>���W�K�x�Mb?�o���ݨ�0*CG����D�7>�U �w�a&�%��67�\�}*���<\�3� �\E�]�|�fcF嗏c �"�/-̅��
dj�J�#,b^ө�)E�Άhk�&LɗF i%<�.�l0]���H�4ۄ� -�#�G;���2�]c'71�&�-)�"��y0C6x�r�O%M=wU8 @5��&^��)-�扽��a������3�����)��V�������ӛ���N�@22j�6F����R|Y����?�r��׶��'nx���Sd�˰$��
֘�+��(E^�wӈ �k���ax�yL�d`��F��5kһ��jσ�o�E�C��6�����K���#w]M{�.��v<�k�� - $��^�INE�	��-+FV�L|w5P0�H�w��4Y~R7��{&m�����^�&�I�-�` ��Ċ�}�n��ʎS�n�$Tlyh˼�!>-�ؗ �j���H��k ���ٵa<n��d�I$�ҝ=��r�"�j<4G��x�N���^y�ޒ�!1��a�Y;�C��^�hy5�����IL�=�a�FW\�?>y�T��V���|
�)ԹpX��zp��`�u���u>�pZV��^��p
�Ɋ;�l������i���&"��]5΁���~q��v���`B���C��F3���YE#S�è��	���g�>�ؗ��� r�~�k������S7�%�'�L��^�:p�3�6�Qp]�),�ǟp��*m�Ya������&y�S�+�)0x�)�ߗ��_Y�#��N�6�;%C���RK�QŽ޺�[�ܓN���e#3@ �wdv��1c�p��ٕ���b�,	Y}	�2������4 ��[��ÄѶJ�?>y�+{�_����aE u�fθ�T6�F�o��<����3�������Y+Z ���.���:��YVLp�qH��q�_����ꖓ�>"O��72��m`����H��lu�J���Qo����n�)e�����$�`;��<T�=��&j�Y9{�%��s����$~�>:��q��=�^�;����'��q[��k0kv��S����,�"hU��M��.�b�AR�l�<iWh�}�I�$"�<�'�:��@��<"LJRT w޼��2~��+sg8��Gw^�d�1�Fǐ���Z��1�HP�薘l�e�Z������hS���7 r��BP�k�[�� /WR����ʻ+AG��Jm�|v�W��L]���@�F� ���+z��w»ŉ9�'�	�=�Bp��X�A�-�y��S��(�8��ӊND_?N�X�	!G��!�y��U��V!�@�����]�]FFm�j~+'F*���{�����U7@Ϟ6 [�E$�\���=6r�݌H9P�G͊j�#tU�A�5�Ǐ���f(~Ki�Һ��"oM�%Vm٨��ئ�TB���X�NG��c���jl�ަE��_��S�5�!1�SUt�#b��� �� 2�s�������_���u�*��}m%��Jڪ����x�3@n�5QSi1-Y��W)	���"eb �ZO���׆���{�8o;)��д���ۇ��jj���{B0d0����V�e��P:,>������q .����y��'b=J�?��i�$z(���jQ0�D>@M}E�x�v���-*f�ò�-�m�IX%u�$n2�y$��*b����\<��Ax���|�>o�!�-�F��v�m�ǂ��3-����Y+�0�D�����Mvv2�LNG���^�nמ��Έ�	��9���U��C�JN��Tg"¶��v���s��M ~U^|�Cw�o?�zt |L�{ꀀܹ��f����Moo������rH�^���
Mx�a��4����V*�
�2ܱ���|���#u$9�âD�@!� ��YE��7̽���އe.08\��PnZي���VѴu(���UF��Ш0�(e�J����>Φ�^�)�etP)�_s4�|�@ ��?�c�m)���!�
��ZXQ&��q�}�)B�_������*�<>2�|n��&�N*��V{��6͵��X��%�����^KtРTȴ�~�1�R�	�����3[0dN��Dwz8"{
w1?ZQ��#:����;b��C���� ��;�	�5��8�����gMB/&�Ut���3���P!L�%%9�Z�(8�C���&������Jf��jV�xlf��A�J�_�^X~Uߪ����9�Ձ�����)�$�)��˃?��z*��\'��oq2��=��<شVJ:�s���ut�;�+��|m��*Oܫ����0�}pe$;��ψ�:���#_��	0{����i�����w����}�9��$t#�N��@�S���Z�D9�r���'�V�.y�^�r���ܬ�|1���_ʕ�nI��K�tG�"�	�&Cx쥵SG[i�͠Z-�0�m�P�m�w�?qɹ��=h�_Ҵ��Z����uD^H�:o	g�P�W�dR^c�O����M�Z�)�����R	�?*¶8�3��Z�Md��{���k����طB�su[ϻ9��h9�%Cp�w7>u��*��ϱ��e=/��91���M��	D�/鳓��>~�a���}kI�S�}Jpg��p7�`A������EY���Bn=�� ;B]%1,��>���B�\���eM��/d��-�t_�m�QT[t=�Ƒeic�;�O�� >��vYWʁX��Y �%�"�d ��.�nf8~$�s���êÎe�dCo��D�!�W�~l@��Ǽ����&i�;.�|�;/���Rh+�ݔ�uWT��6׸�q���D�#s�t�b�6j�t ����)���6{���
�:E��ܙX��J<�7��n�$������zlS/���#�84;zG��Ň����B٪xUP0U�{>��R{|�@�v��["�K�k��A�$��G_�A�hj����\�ie>�1
���؍���Xݗ��9�H���W�-���.J#�wu����2��R�gM��>f��?�T*������Ҿ��S/�'��3\M&�of\��·��x��D����ɿ��e��\�9�r�� T�,���f�J�\kS��5�W��k6-���[�zy�Rs�U�d�H�S�4��qK�pu������m��],�GcF��W_@��i@A���X��M������wlM1S4�FA�Mc��7�~S}�	CG���\��8]`�-��^�)���YJ�(�>4��ǅ�4� ��������6C���"$LN96�kӢ��S�������K���oދ�4?b!�=t�S"!�srsg�l�̿$��ye��9AP>ڸ�4���/����^vy�<~;fyi���,p�kɚX|ȫ���'��V}�`��&e_w���c����a�;a�1�ܜz.���
���AP���d�ǧeH�6[��GAZ��ӭ|#p�ui�Cy�Z��,�$+3� ���R[z��� v|�u��G-sz#,��yݰ ������)�xZ�3*�� 5B808�r���%Qx�ܮ�#KѪ��9�)O�pb�_��:��W��$<�d��h�E��./��$a�,�pnW�d-�%�Ѭ��>��ƭ��~�̻���c��ƺ�x�+����b��&'�4�E��Ž�?o�6�Y��FE��w�pw;bon6���F�ܣ��8�r��z#跗.Ta���� z�a�1�v�7V�����`�$�G[Of�d-���,h���ݑ6z��T;a����"���9��cM�� W�U��}�����_"�Oe��y/0��9�v�gU��	ʗB�I�Bug)Rʋ�3���$K(�@0�:`���/���r'�rV�<>B��e:�ץ���X9o��&j�o���Y��4��>��iZ�R	X��X�[�Cǭ6��#�C}	�V��^�y���E��ͳ#~��W����ݱ�Z���DN��Fg(��l��G�����R�_�Q��RԷ��5Z=��f6�b����㥞���y����w�ֱ�u�PBV���T���B��1��A�"��U�Z����@镥�B6Wr�Ƥ��
<;�?YX��g$Y���7ʁd�1�O�d�O`���-�v��L���FƉ΄&�ޥ�>��#{k,�[���f;�Q�Zt�0D$7�PB}H}Q�925s�65�B�9r���Fe/j%X���A�q��>N�~��mQ�sl=�����S���؉\z���@*eM'�$�Λ9�?�Ia'np��9pQ6��׳E���§i�
�"0��@�.yJ��TTjM��F���X�}{�;���]F����1��u1�͒pv�&��47�K�K#���6?��.!#�2k�D�-"���>%������,�&+�P|_�ȇ�|'�x��6g/O���6"P�B�������gN�<�{��x5u�ϭ�f����{A��2"���r�?�3ޚ>��\8D���OW�\ 3-,�n8�l��0A0���xZ����ԏ��QCdo;SC:�"�y�]�cD���QH���x�>�@���.�giC��۽��+�F��R�?��ν.��N���6�ϟ�|�"���^�(�X�>��b�@�b*Q	��
r~��"Z!��k-�_3,�"rk�-N���m·�+��D!cV��f귳�8����xL�7Dq#����S���h��[�j9�`��ce��W�8B�4��ćý���,�s����8��4B������OIE�K۫��}N�ǘ����Q���2�E��f�j�V���J�b��'F�7�^%�wi�=��X?~.� nDL�/��7��r�6��7��np�o�f19�ǿ0�0�_�Ik�O�͌�����I'��6���9�1�Vئ���ݑ����C�YH��'l�Mȹ��퇲��8	�2:�&�sԨ
}*��)wm���5���n@�U�(I�/hZa5UX�C���ĢC�Y�	W��;2��Ev7Q�c��������Sh���(�:J'
]�G��[F[jiْ�?�`zh�R��O�g�a���˺+�n�>�;��᭕�f{�a���������:Y?�(�~�
s�ԁ��#��q�g��&�z?fu����*���z+eI7��!�B�0�cph����(��c����>����`t�{��ԱFD��֜�2���
�tx]�5�~Qm�m���a��?K���s\��ݿ~|�e9IxLV��I�~��D���	��ߗR4t@��l��J�G������ThS��\8�\v�?l���/��x@~���Y�0T}�SZ��|g��n�2^�hp�{K�6�O���P�5�iAVp��O�M�k�����1i����W���C�tS�r\��S��&z�H��^ـ-�>b��?@�v�uq�훞�4Y����{vƻ�R�����V"q���όr=F
��,�[o[�R�*��H҃2�m��V.�cLͷ�^c�F��g�P9��Fɛ���qH� Й)Ţ~z�r�е�`�F\��ݚ-��K��,* y�EvbtZL#�%���X�����ZzT0�F���A��l��R�S�BLp��� ��@9�j�y��T�2�`��q<;.���>�����ֆU���/\�Wj�/�R%8{�י'��2ǣN]B���UU8�dEp�r�Ǎͧ�Ҝ��(8��l����NK=L	2����z�d��4ͯ~Q����AI�e*[B��?+9��EXN�P\eN�؞L{��#� ߤ��ƻ	��P�j=���!e�#���BG�ۀ"+��)��N��3�OV�%vA.v$*��A{���lt�$��q��.���@����8w��+E�(���J9�s��>����� w�W�m��+������.]s��=4����#/���
����s�۝�:��?^��#*��S�G��r�ka��y�?>�ӤF�+o�U6�c(�Z���)jҏ����F����8�%W�@A���w��w`��<����0�C��,���h�6�C�R<�ӃU�R2���e_RДHg7�
�9���
�n?�i�>bLje#TU;t�(b�~D*
�)�o��\�;�1B&Q\9�t�̔��i1�.�B[I��k6��-���p�[z���ȕ��Z�?�Ց-���| �+��Кт���P�'����$�������pd���7�3W�u�ɼ��ELDx��?�ر�p���Q�5n5�~���C[R1�{�[�X�6�+�q1�*Ǝ!%܅�j_>��{ը�7��K�zx5v���
 ��U�[;璛"�bY��a&����D���3��5jlZ$@R������6E"�d�Vb��N�i=���f@Of�H����S��Ns����>�m40PDz��:]	���"��SOK>��&wVH}�~���;��6\��Y�����<��b���[ꂸ��=:<I�_��x�����a�d���)�q!����^0$f������`�b w@�h������?~]�Z�Osf^�Kd"��/�gM/�����-��j^�Ժ�ױlH�Z"�" �]t��#�Μ'x�o�;БưߖŻ�,���e��
м:	�[��g�o�������&������+�g��/47���W#���-�(Y���J�ͩ�@����isʢ�*�dv""���=����ˬ?ɔԊ+��x�q�-����q�cG�@oVK��P:.�rB�}�pN�BUBM����Z�[*^�yo��#훭��!��d��k�>���Bɿp��BM1�E3#7#r��
����OFR+��7uϭ偲�|#bda�}�~ӉCX"9�����K�=����\�_fX�K?�Ba(�_�Y��g��0(���t�t�[�G����r�y� �$.�m?�rs��/9���j�"*_J�l3(y�<?���ȝaC$�B#͟�N�`�����ěL>��|�.7l1F�F����ާ�w�~����!%��^�Ov�M�L��C�@���� D�I�>8Z����T�0������ٝ9���ت��U9��Dt�:�Y��2ʵw�T2�,�	_|��r^���C�`���1<�,t*'�z�K@�y�*�9�X��c�j��=���Rm�3��9��̈��T�M�{l'�C8��I�ťe�4�Pv[c��d�����n��4̳���bf��3f��ϼ����1�v���7#(9���������#��h�N�� �fH��7�=c�0�/���y��a��̣5؆�����Lc9{c���k�CF{���́-K�J
���C���Hͨ(��ғ�a�Ɵ�$(�0t�3��XY-W�fV[��Z�����y�34H8��i�k� ��k_����h��E�=� �訮�'["���^��ӗD�����9c���H+|�q'�}�B��&|���ѻ�9EbǸ\�8.��FjиT��&tf�
ݼ`�iu&,6��>��*>�W�|�we^���Y-FW�.`��g u��o���#���}�����8�^��+�Cd������K�Z<R���B�~�W=;��N����t!�v;$k��F���}X*�RKd�������Y�zɕ7xҸn.t��v���i�D{s�V��n�5��k9S`�����:�H�jT�{}���Ò;Z�à'ƫ�>��6��T�\+���-�j�6kݥ�>5�$��t��?d	��"�U�����	1M�O'�.x,:]dD�� U�����y��@��M��:�7n�Ϫ&bn%�3�������t�MT���g#�N]s��<Ƌ&Խ��Mr;;���m���ľ�8Wa=�*Vy�9��{$2p�{�;U��:B��:q vB�3Ip�gt�D��Rŭ�$Y�h��n�|T&�^��I�5r.������#�o�A'��ir5F(*=�*MV���d�P���.�3��+B�|J�ˈ�O7)���n��X6	T����C%�l�b���z~>�hb�.S� �y5� �����L���;ތ���Y�v8Y��'��-:d^���p���͕^v��Y`�\��lk���c|�{!������]�8�l���!�+c���Ęn�/^,�fOܽ$m{��0� R=�Я{�[�x�J����e�~��_�X����2���P��*w��\���V�@���jo��9�?��^�.�Ot^�T�|�ѵ����2�я�u��<#�Wo���,��R0�7���Ii�`�[�		�ĭz��1���wr��g��:�=�js��;f�F�u��8�2��H��jΖ�����[��,�������l���@��yZ<+Η��F�l�\����tj�>���V;�KJ+)�.֏�V~t~|rc���BK���3�4~
���S�g�u$>uP�)	Ֆ�������C�_HA�]e��6��Blun�� �v�- ��".#$�!h�����Oz
@���/(�P�('c��>�<��f5}����]���>Z�2I!Rx"����)\�ח���0Zi��E��А�BW�t�-�&�i�p�KGa�pBO�l=�L,H,ե���Wj=&�����9XrF�n�9���o��:&���W$z_t��6{��n
�U�d�r��a�/��U����$\׉tk�cf������_(;`]�V��_�HP����X�n؁�N��.����y�~Q�{cqz��O�$[���:[ɿm������yg���ÜE-�i4�V�˸(�0kQ��%��;�s���A�&����X�0bV�@�4W�Ub0����<�.���r�P��Y]TSW��fΰ�I��`̼����r�AeI֊	��syV��s`���Y�agnl�	��6�����,��bC�<Ҏ�r�Ё�� ����>��D�եMN=s��N��S�}W�((�)�0�i��_g¬1u#&]G��FYSz&��0� E8���nB��{f1�"��`PO9�I��g0	�^I�������$��O�f�E�t��Z���r�b�n�p��Z����H�1
�s=��%����`�5���sTj�{n�޴K⸇��.���v�����}`�BH ����8�$����?C$f��o�0�]_<�D��$�զ_�}h���~��>���o�zIv����gf} 'Ϻ���I��,��eN��'� }N�5)&����UmqLsv���hoϏ�[~��?�$�g2^����v�îA��f~
Nqa�<By�5��C��|D�,�VB*&�-gQQ�kyE�������ڹ�SҔ�l���F�n�NB����n��H�w��{V!���D���@E�q�~����U^�4Y��C^�+��)]!����R