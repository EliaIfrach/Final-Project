��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��-�ro��i�����/L-�U��lOjj�l]I߫�p3^������_"�'j�ʬn�*W�� �a��;��}���������)t�X�|�r|�~U���;��k��2��%�`�	�c͜��d����/�OB��*$�K�[�>�)v���������~$�sF�]����ZP�6͝*����ĩ�';ɒr����YU�|��#��Yq���65��~�Mduث6z\j���4���E_w3�Cن̷����o�I��Ƃ�G���~T�VO|�θ.YW�9�����I�0�J����r�=fw 	`2K�$]�NF^-F{Ux��L.2OP&~����k2���S�BY�F���iG�H�E��+�%h�<����I�[��G/*/�F��➳��nZ�W����Y�o~r��_�$��\����f�M8D�o�OO���"��D�_U�@��MC�`��.4W��ف�O(��
��,-�h��jn<;���#��'>�鑩�!i����8�1	ZB4J�yY����p>G�����ٯ�`����?C��?��=Y%!��b�IWx+����Q�XjD�I��5��� \�u�u�@n�X�gs"ݚ�i\�X�8�xt���'� �� ��\U,��P>�Q}�������g�]�JJM,��𺪆l�
��z�G�+�QeE"�<���?�PS��"V������FSh�Q��p!�o���M|ln�P2଑��\v����7��e5h����p�C�M"�-�v��4͵ȁF[�=0�$^��ܜ���y��Q$u$���6d�
��"Ｚ#�/��/���34�}��$3#|���2���"�f�4!��Bˢ�mn@��Q!5���SU=��h��qJMr8�q�<l)�Y��Ѐ��������eg�fMV��I-iҷ~$���^e%�����^?⬄�٫%����@(GI��}],#&�M��Q�_�z�-�e�_ ��Ԛ%yQ�?��ǆ�3,l�?�|~'��m��2:��'�(Z;��3�bW�O�w����	'J����`W4xx��Z�4��g�d�YSDņ�y��"o����cWHQw�y���!�{Q�����6�����]�������oh�+`A���i�+)�(�h��l#:�x\�9��J��HϽ�gx�\�s���j�nc��kߴ'
���L^�l��r�	+f��AU�S�DG-ң/�]�͞`5Q���X�խ?�C��;z�Z*UC��e���ď���?DzcC�;ᨇ3�xR1��J��=f��#����+ *hx�i�8�κM�$���\����@֝[v�������r�b��h�z
3�jMlK�U��7���q$�L���J�'�6=�
��۫g#�!���u���EB�Ӳ�-��ۮ4�n��V���	�(�K���}�����s� �����*8why"��6��Nhr^b������@�pGD|	`V���9�^$��|E(�������Z;��p�L�׆�M��C�Wi�  D��x8$ӹ5FW����ڞ�h�"����,�]��tX�a}u��{V��wm����$��
?��7W��qlI�L�L3���O�y����j�	̄����#*K�8.�'B�^�ؾ���h��Tt�+��}�"� ��؇��g��~y��}�K����G���M��a�UG	n�ݥ�%c&#���l-@5��nD���8.�O2���@b��-H.���������:\c�zf|^��F���za|O,�r��)�i�?�4�ln׽��Y��
< _�km&�=S�0��"p���B��z��"#Bxf����}�J��ϐ��i��G�|R���ӵ��Y!���-lT�t��ӵ�T�Q�u�&i-ņ�+Jw"{�T*���R6Cz��Gh�NG�������
�(w"O��'�&���I���ˡ)dGl�/��&a�:��vU�!��L9^v*�w���;?�������4�tZ�!T�z�X���Nlu1)W�l#�:7m2���׈#s�9��{�[��F��"��e���A�E��@��j�˴��r�l Nd+.�ǰ�x�� ��q5A�0�/�ٱ^����1g"g�au�ǩ�9Q8��u��MV�I�����˱�� �LK�~3�^���)W���E'��=7��N]�^�����P~^�i7��iPƤz_^����C��L��o:������e�ER�	� �]v.9l~ۇ⮙yܕ��>�R\���^�}[�'�#l&��r�U�i�Ԇ'��r0e ���LLąe�\��{�Th��#����1����Y������Z�J��f�6�&�g�_�A�6��E�T��4���G2e��\Ƨ;�}�QZR'�6J�d���¬Nں^-�sgS�i\��`ێB*,>��r���Ҥ�Z(R�;��:��A
�B��;���mǝ̶�c��H�����nY�N��ȉ-wg8��Tu�9Df>%�in��m���o:��y�t'M#߲W�1��g�I�Hxmy�4�M�v}���-�C���|�^���CJ|Z���T4s�n^������R��=>���b�t�H�|$ĳ��p��d!1i~�*~�a<�:)�}*�4�����m4iV�+���o�Ÿ@Sݍ=p��m<A�0��
=p����+R�=�2E�bzq���u�$Ƒ�]4���l��¯�q�pqh��ɔ��{_�y&#n�Y�? �/݆�x �0�CvO,g�Z��f:r���Bv�[`������\d>A;�=2\6]��p�P ��0I������{�B``��^��U��O���~�]�x,���������l�j���>��*h`X�����ݕp!!@��O�� K��)��jv��ʦ��1��cɹ���N�#�m�j_Æj��+�mK4���'�.+�uj���en���v��ώ±�@펐�ݶR��ss#:��X}q��8d���q���?��{�5��3f���{sc9U�:
P����s�0?���Et���/�I��k��{(�5yL�'��ҋ�aN��.�+�&��×���Y%�~,Bx+s�9�LK^��(;�Q�a��
�����M��ئ��d�#��3Io�-\�
�@��eAH���B���R.�^�z��M9Cp9%�7�/�Ǚ�ԥ/ծ�Y̖�e}���֊Y�m&x�?
���~Ӡ��WmnFs��\�5����&e���GRĩ\���S�����f�G/��8*3T<x|�c~�q��W2�I.� ��t·��2�)X�%@B��z�����ً_��L�@��N��m^o	��mT�ⲛE�{���������d��>�ó���֠��;�c�: �`3��f8�$�t�/�͕�FE�˗
��>
�^<��I,��@UA�ȕcx���z ��*�)���
GÆk.s6KS��
)��&`�v]�oӂ�MG`����BP _"�7�×�5�xR~+�&~
t)%�-���?K3i
�xE�_���.�o�^i�J��v7� j�UL%���A^=?Y�·I4���"�°g�~���.�2�x�]��
��s�>d"�`$q�M���T��a�ֳe5����`4\a��Sn�G&4Nx���@�����΂!�3�>��F��Ua_cF&��~\�f���o��).k�Ӫk�_�4���	�M¡|���_/6���<��6ڥ�PFD��&C�0%X-�h�zb��!�qc���S����"Z3;\�=��{�Z����3�R�#���V69�H�-�C��1� �=����fs���,hPi�+�V�f�ri�8M���H:�*�5����C��t&l�}�^��iB+�a= ������yH������?�(f���]�v��'�̣jNY��%�'f0n����������w-��Ͼb��y��!�x�܇>���1�9x|$�.S}��� (V�����N؈W��dTI�
�)��� W�B��zp����dY�{�/�p����L�J\���7S� ��V���<Mt���� h��?�Ck,?}%�ư]����Zw ��:o'b?RZ[㎗���x����%Ň�����»���-��u]Af��ܽ�R��h�BÁ�N;�b)�|���;��}� \��y  ��st�_�+�obѯ%A;�[X�Ԋ��: �����y�-=y<��x�+J��~���ئ�O� `A���1q�3i��5�/Ȓd��w38H�KX׿=�s������g�Ͱl�۩&�5��뱌*Sj������s?XB��Xm��a���EG�7t8���gPC���5�X�
����>D}�|�:nL0�_~�� �,Ɲ~dKEw�F� Ak�1Bʉ��8�KV�d��	zN����X�!�ͪ+�T��J7,�~F�V��Q��z�2Ͼ��S�z�I�c����?4(�L�������Pabw6�I��CFtt\�>�����b<=����/����Cz��8"�0����h?%��,�j�k"��m�ZL��d�%�"���7��ː�����E.�ɍbEN���S� �&��9�D�6���N���:�|m�,����)G�RQ�D�")�!�S�X�n�7��Y��TN�3&���4~���Z���
	)�to[�i�����1D��f����0G���F����q�\ʨ�IOݜ5�k˻��b���Z�� �X���J$c��g7���݂���