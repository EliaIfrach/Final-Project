��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
O���w3�?�>���*d0�vjq`U�ekOF@6.ђ�ᣅ�7Q��`2q���IV���*>��N1����El)^�&�l �s������!8�(^Q>I�!�������a�bmWD����!ut��n��]�p�?bk�C�S>��Yb`���y��є���M6��=8����۔J�0�%�G}�1�R���	Ԑ\��p���;�?��o�`n��7�z�藀�>nB�ػ+$y����0\{O���S���ft�9�7���(�ǰ��(3��~ �xvfp{�Wmm��)���)^�*5H�<������@r-��B2�9{�̽N @^�����_����\�����A�������'&s�����b��S.�x\��.?���we�q����7�-�;��԰O�#���)y�͸���w 3D��|�=3O9'�憩n��)����.vG�a��|\*4j�k�x��:�5��2ǅ�0[��ep����K�ֶ���	"�,�n�X��ڄj?oK����;9��{��qe�;#y�6�K{3�w2�$d���I�V4d"#ƌĒ`p��^�9�;A���J!�0�F୨�Ռ1�U\�jE-S��%���U��_�d[{�-��_F�K��x���㫀�Q�&}�vh�Sb�b����:f�J5y�f��m��o�d��*tV��'�����4���Y!�s���5�l �}��jY.@_�ٝ7k��{�/�앿���Q���_�.R�%g��D�'�:���j�O��n��nLUD(|'V����0�_���a2�Hs�����,~��H�|T��D�{-�*KvN��}�<|������n�ڼCV���-�;*�(����<�sz"��58���OTv~C�|�!\i$��Q�yHA�y��2��]�b���yL��I��Wpڟ&��k8[��GҝcX�͐�>}�=�Ō�*Q�&�!�$��!����Ҳ2��꘤�Q�$��rB���K�I�r�T����9)��#����/?#�gU���W$z�O?X
�'����o�2_HEg�b�'���?9]_��n�b���A@�T�r^6� | �䗛�7_�]	���L�(7;R����\��	�l��8���}��8�W�(�^�R���싕��n��w�� ����e8sb!,ێ9g�ʿNL*�n*�R�sN�!�X/zTH�8>4�i�XRλE@�щ��������iJ��`��T�L�IO!��!n~��*���������JD��\��5��,qT|�3�u���^-H�CB���&ȓ�C�#�{?���ݽ��ck�\��
�J�'���J�<�;)\�6�1=z��-���`#��d��g�/I�W`��//��W��62l*���B7l[��g���2��7	��r?�`����/�T_����0�=��Q�_��U�d��_ө㱶��g��if����^��hCl��n��L($;�*m��Q�;���&?u��h���1j�@f��j^{�@���]���7�)B���<�b<oɚf��=R&����"<u8yX�) �G_����U_*�, ��Fx�Q�
UA�j s����ȳ�g�Ɛ
�,��/0�F�'�O�݀瘄�5�i^;������>v����T���Uz�H�W'�a0sJqi���� �L�s
q 64X�i�C+fTn{���눞'��������E�#���|�<�sJ�d�N��>�{�����e��i[��1n��!�B#g���P|��>�J5���,��+&�|��}�?����7�(�23h��\B�K�\U���A�Žum�a�4p-������vtA�U6E�i/���0����X{1���I��da|9I��=�}Wؤ��4�wƏ^<��?T05�L�b��3Rmt8��0�#����iFC��{u�_ݎ���&��!Fb���S���3�.��D6z��[ċZx�ҩ�)\7ʄJ[?���ι�{A|���L��a�<��F�YY������,�8�H�}Y�ʭ�����KX"n������=�bOܶ�Ziɟ��Ů��X8p 8�#��l�}���Ive]���̾G]cq��vX���'!�+�����8a�"r����XfA;�'�zo��#���}�(Nʻ�E�?���K��g2lB�NzMQ%���ލ�{#��y��aã]A�yH�醉�ń*>9��CP4esb����7P<��jbK;��#ft4=�ߕ�.e����A|���10�/�E:hY.&�y�DKe��5�u���i�H|�]�$�NV3)��Ҋ��%A�h	PG ��HW��皖k�Wa���U:ꀦ��j�10(����Pܻo��%��\VO
;�]U�H�Yx��7C����.8�$��:��}���w�A�+��4W����I����i�m9egiJ��V�ґT����u�/D��b�����=��U%���7H�o`��(�?�,��Y0��k�������,`�7��A0N��#��O]�A�-N�`tߒ1`�/L?�1�{��o����7 i3��s
cI_+O���A1͝ %bʢ-u�q'�<�n`�j+��g
��?�|��KC���<�9�n�	��8mӌ'阵(�o��.f��P��	oodA똍q�W��)3�:��R{e?G���ë�"�˩����'�u�rr�ZWR�nGp;�@I^�ܣk�S��zi{NM���=۩6����aʆ/X�ٷ��!�,w�JF���3���E�� ��/�=�wC��#7P�x�����}ݴ`M���'X�LPP��8�|��\��=��惽oO_��^`�ѣ	��� �27������<��~�L��rgO�.KH�cφ��Zb�c^��>�����{�|l�;����n��Zj�&��/��4:_w�d�['����(�.�$
��3�+�I����<�[i� 8$���9}�&sA�c�(�X�2�lɒE�����K�>�LT!�n�i�ڱz)uV��q�r� ���s��gPbH7�!�]l�Z��_<��qa����(@��NR}O
u�_d�R���0�/�~F�dO�=�fJ@|PٴM@����X F�MR�-Ⱥ6��43^+������D'�4lČ03�K';����������3��\�fXHן�?��@�Z#��խg
VE�����q�\U]4��@+Q2e��hq��+7M�ä��Rk�wo{�d�������Db�2%������+���K��T�>��� E���
�"��Z�q��7&�����*>�L���.�ϣ]�y��IH�$���Ұ��r�)=r���h/MR��fߝ����P{ Q����)��]�=���IYdu��D����Ѵ��^>� 4��m(M̲�|!�҇�pb�hv�{���q�|���^̓�_��)�u�q�]����S�.�5�
C3ߪn[K$�=���Q��Uh�����h�h�����*��~"�Lʭ�$�@�=��Ίs�¸ѻG ����!���1yV_����(kn>D�	�]4? A�A���C�����
ε��&kQ��(��: �:�̎�ap�,@�C�3[�2 l��I�Ӈ�B&2�;g��7PkŠ�pm��cRD=��F�-����@�,q(�V���j���Ju7B� >�فϦ��=e�A����6d��@�6��">Zs^��k����q_Q{%)g-DE�`�cUX�a�./����ojٕr�K=(9�1ߨ����*g�P�
��=�)J̃�-H�v'���瑉�p,~��x��T$�L{8<�$3-�䊾�>з|LR���h�z5�k/��������6Z� \xR$�>��7ں9D���jS�4��0���G��R3 L�#0�{!]�#Z"���S�o�H�H�n�Gˆ��_}�r��iު��9O&�40U ����.\��%r���uAI��hJ��ǖ���q��r|�W|V�Z�"Y�!���	w{�"rSY�&��QcŮ�9sH[s{C��(���+&�KOo�A���1Nc�u��e��?j��y�Ɉ,-�mW;ڐ ��MXOtK6Պ�3P�ѣ���ڍG+��9_�<J:T��Z��:��]%ᕍ�9Cn'��s�2U�ܯ�Y�w1��(��%p�e�Ds�������o�t����nkG��*���_ad g��@�n��m}S�Q<'O�_iʔ3�
�fY$m�=��:�f�d�=��fK���>���͟��YH���ϐFt�����hO.1�,a`(d(��!�;�6�l*&��d^P�h����KR	1����ݟ�FT7N^������J���Z�O�����c�p�A��F���ˆ���l?G��K���e���_���8�eo�P�<v��-NLw-��U}�w�֎p�v_��ʂ=M��.7��t�W�{����l�m����x���׶gA�����K2�L�\ea�PTO�/�q�ܐ����y4��	>(�RA'�tu���ؓh:Љx�P(�|M�I�fj笅�d�S:*⠘��������e�x����:H���&w�|W�0�?Ef�c��?x�Cq_�;�w���)%90�+}��K���y֍�"�Q\�7�n�#Ӯ7O�	��R���R^^9�)2�6��S��gMލ�l�I��%���&��d%	�,��f[�м$��A�(��GuH��6������s�٠3Mk��p���M�Lm3��>��[k�b�b�����7V�H˕n%��S�V������py�ؼ���º����`�Z�G��G)�%4���t�!,�@�¼�S@���u��u�-�(�M���\ŗ�S�t�PŽ"�c���;��t�6+��5�`mK2Ad ���t@S�Ц[�G�Ǿ�铀<7q�OMQ����vX�#�vP��bق�lu&�
&��gi��q���Ռ툌i'd%�l��0�`�kz'"��Ɗ��1J���|	�rSI)�Ū����� SG|�fº?HS!vn�b����f�Qu2����e�mF,��Pal[E��H�q\�LU�e�,�ŘO�9@�m��@�fc%�����M�j�.?��<���.�3՚��A@%3���������5�d}�7ܓnV�b`�,i�+�4Us�3	dC^��g�K�����V}�!������٤�-"��\=F�w`�Fh���\X��לJ������?Jfi/�6�q;�1��I�`�h�N�;����uJ?}�~W#�n��