��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
��e�����&�F��fu�O5?N�Oѳ X^��Qٱ��%��R+z,fW���;������\g�JM�L�$�B�}��UF�������7ks{t���RFq��j�ȋz�n}*Ć�/�����Q&ʶ]Z�z�=�_H�������'�&���-4�=o��Iag=���n�^1rչ>0�c�F�>�z��8�֒]���b>H4(���]	������]�73��YCr�񱱮��PX��K���(O��2`z��"q�p8� ��'���]u�!a{C�F?EWq�b�a8x���+�H2�rX]R��(@�v�M�Jsá=��o��j���괾C{gX9����;��A��8�y,�a׬���V�LDѢ������V��E���ŗOwX��ݸ-����ͬ��\�;�u!��Ԛsg���t��+�x)(��Y�nxC1��ɉ�~*9�*?_�3�kL;��T# vP<�{���z�.>q���2��ǚ0@����|��?,��+�˞�ś�i�z[}�ń���!�!�)尟�4"�٧2�)"1v9�+F$�|�f=x�aD���%^�g˩��ڤ�JT�7
�lo$y��U��l��Y&y�+�E��K?�'h�7#J�~��G~�g�TO]���H:����O���,�X��+�%�c�ܝ
E2E��
�VC���)�;潔i(ﷀmp���Xf�+�['�)�T�M�{0�+��v� �(�+�[�~`eءf����b��Տyu�	fL疩�at&���9Ƥ��"�w��C��=����m�/>�ӝ��ڔhv���.>c��	�-�Is0^c�����u��u��P>~��d�N=p�S׵59M���$HgO|�fS���λ�~�^���D��_��9|0MrN��!�ɻ�3<�6)�=��מ��O�W⡅.*4��H@��9X��N@���q)�@uc��!�Cv�tBQ�Cv5�p '�ߛ���W�#�v٢��}�:�/���P�뉶�SBU�_�R�W!�����I�R����t��.	!�B��d�K�E����o)���Z�&�ր�;�Dp>i�!W�Zh�dh���5��R��d����j�Q�4\cg>�D�n��&�R�߂n���'
��S���@e8��ml�/:ȸ<?+>�OO���,�_d�Ҕ7 -&��;�aЅU�b?��YR����șRl;Q�0\�(��!�v\��ᆛ�*WV��c7x���}�[�������M8�,��S*�f��7�Qw��ql����ja^�鴭��_�.0wZ�Z�s$
���s5������M��ncYK�k�m􍈵U��f&�{o�_�u>V��6��ۂ�}j���3�-R�ވ��Z�Y��8�t��rF���o�^p�\��Je"�l@�R|��ER�O՟+qqd��[�i��d���W�g��I�R�p��8�RiBgfϷ�M�f�[�Q2:�}�4Zrc�}!�γ��U���"c[��:Y{�F���C��L�\���aH���zq��r���`S]O�8�VZ�ׄ�`ys�@�;F������g���ī��tyD	`�[�jD�-��4:��fp��]%�=�TW�
8�\W��

�F��|�:oD�%����w�]I���U^v���^�5� �ZZ�-�gr�H������Bs��G��/*(���/��_A��{�_�����|@�s�*���X�N�n�giGo0�>�����D�@���ߘ��oC��2dmX�i09n
�K2*=�7A��:,�2�ǮI���A�hL(���Wo����#u���6��
�D��[��9B39�𘁱���Ҥ�|��?�s��/(�gX}׸�H�P�]e;q�U2a���{��F�x��#gh�(o��{�h�����v�B f�����|���c���ze�F�H=��,��������������+[>ج���ZM�R&4�_��;~��\f;��xN>	)����D\�w�ð��JY���4�7v��EAXAФ2��N�����O�8�t����Y8�o�;����+��ZƠ�M�A,��~���������~�}uTS�1-T_��6h�9$>�NX(�Q��=[�MF���7���vb��| ����s��vK�@:Aj�)C�4Z��c��F�.t1a���;�AW�L��,��x�*r��~��x>���׵�J/� xw�TW�v[a�>6V:_�L�-U�cJ">f�F�����1û��0@�vԈ5����2��T�pl�߳K9��RB��rz�!u�^��\�fB� ��^d�������i<��ӯ�}(�'�z�u��8�Y��	;�Ct��7��N�A}0y&�� �Iο�9�I���;?����kc������G>j����Q�(W�O^+G���� ��F&�t寷�3��  X�Wc���N���֐�8����Y�l"2cZ
�I����uz��U�7��#3f��?NE�.S@�=4:�v�/�g�6�������[J�}��
ɁN'.e��f<LNb��Jb�F1��,�k��8�"���![�l��?B�nv�~a,��	��}��гt�p�.�E��C�,_w�"���\1�J�{�YJkEոUU��ii�A��*�����MĐMW?{uz�o����en%zҗ/eC���m��ؤא�EI�Z�f�%.��V���i�����K��;��u'q�D)�ۀT���DpQַ������JxG�G��e	(������+L�$H��ܝ�v���5_��q�`b/�Y&ʓF���^��7����f?Q�ې�fC�;}h{����A�ʫ}0�4��ݚ�������+oM��o0�V1�]ZvH�_�z�S����Vǹ`�O+��9KcYa�Le��b%�3����W�SU'�! �A�^��~��`�L�`���FR���}��<A2j/l=�o�nD�^�%����V�!g�3��z����{:W2�N>đ� �.K(2`W�9v���7=���6|��ȩ��M�v:n�_��?wap�̳]�E'	����1􂴎����b����O���\�'��%���y}���yJ����	��'^�����+����>�5�N��vKs��������&b�I'Cxk����1L*�
�����;��P;/Y�L�ׅ"b��'�&�A�Ԣq#Ǐ���ǹ�ΜP�B�X=IY�;�߮[W��졭q�~�9%�
;ic$w�7(:&�yx�0�3}�r)(��AVcaM3]z�DNݜ��r`��Z��0S�]�a�D޿o���5н�5 h_�{����q"���|T�������@Lb�>�}�xNaq�AL��śp&��gO7���{��57�� ��x���R����Ԉ`��5�)��JJ�ϗgmΈ,8���N]k�����z0�t�1�	^�6����	׶�����b%�����^:#ᩣZ.��0���F��P�cJ�pO�Ж�����'��0�֯GbO�3���gg%;���c�B�۽�.��n��U�����;M�*z\�܆��0ޟ�ZXB�\ho
q��'�iŔ���'�Щ��ew,�*���h�`D���'���Ѷ�e�,}�LPn��䱁 /*�0�t���L�ģ�-� t����o@�@�_ѴL`I�t{_9A�*���xD��N}��M��m���.��M�3���o���N_�;�ḁ*���p;SX"rz�π.Ѽ*p�:o���qrb���i]���Z�]�'#��4 4S�l��ǴG�Lq�(}�%J�a�W2�����D��a˺z��@{�0c�i���W�����3/$�LL�v���U
H����\���+Ė�ȿ��L�7�'�R=]_[F?��q�(bCj�V{�U���d�Qe�d�_5^���jDS�'3�����*�Śߣ�`E��
S�~�V͜c!UNe�v�e���o���ʋ��.^&*��g ��\lr�n;����~�1܊wf�+��:} ��S��.<Q�q�|Q͡�!���\����i���G���f��JC�����Dj��8��yd�������ڗ����ȇ2� �đ��=Z3�=UV�y�5������CT,`I��l���o�j$"�~�b,�wA�{qp:ɜ���M]((tV2&��)����$.��TxL��~�@o��2N]4�}T�@��)��s��rpPڹ����'�������� 90��������C������[34�(F5T�_:y�4�{G��l"�s||H��&��zxfD
[�u:���qɿc	�o��
q`2��g��ς}^�:p:w���JKU-�@!�"���&��S��� Hce(�M���F�g@w����yY�.�$�R��#ko�J�|B��E!H���W.{�bA ����|��S���B�,��9:��̉R���[;�X���>$G�(d��ݡ�� Ӄ��	(�%���U�o"zśT�L�2U=�=xt����q)���i�h���ЬwW�;��l�Q������V4�*�9:J�+5P#�!	�W��֣ ^e<C�'V�6��v}��d���vTR����:;�&����H
c+�A愧YR��b�gez�%��v1�[moC���u*� 4���S�8�i�����C&���Ib��P�+e�ך�j�Յm ��}֫����l���-%�&3��-�ra8xUl��%�6�m(����;�z��Tځ���Hf�s?_���vz��Ձ9���L�_�C�K�,Ur�#!PF��M��B;�1B��HU��i��]r��8NЫ�^����ʆAf_�5��J�m?����2[�������� I\74%�w��3�ra��p�(���-4�����m�ٶ
�����
X�:A�⢘P�'g�=@�W��<�� 3��q84q(�r�T�ppb�W1{�I����U`8@��� �u�Ԃ�("m����@�`�"������l��ۙL��߅�|1�!XB��Q�ĊC�>��2�(Ë��u{
��!JL �aƀ+�R�{���C���*}/N����! ��	�b�̏dTID�&�^n����^�-���Z�L"YL�X�3��F�|"�A󪡏Ny�D��� 򲨄^f�� �V�ke��
��QAXgJb��>lpK�7���(�G�~�,�����mЇ�Y�12��*��Q�S�E�'��@}��� �%�{���"F�����&f�[�T�?e�ō�\]F�'���fdi)��ͼ5�����M������	ɿ2���	���{�QoLoR�&�d�A��#?��]��@��a��h=j/j�cn��A���=g8��~n#Ñd�(�X�qf�������n���8��KE\�QQ����G}�g&����,���<*R�Z��:�=U�t�ŮbԌ+x�����(���[�0�����1.�m�Ia�S��A�g��Ԧ�b�9w(Ѡ�_uk�?��fj�z�'"��?��b#m����.7����#9%��*%��OQ�D<��ڹ���-�i�@3�{~�`E������?�2���z-l�҆��Wd.~_g�biњ�'�s�<�FC��9<�D�|�wc#vo�W\z�����Y�P�%�]HF�ݶ<�������S������|Fͣ�'�Օ��@����D/Q�Y^�w�s���{aYHTː.�������P�B�~T�>�d-�I��6+iŌY��ߵ3*����\򳩸�	.���.`�jDű�v�NG��� �$��e������?�Bu�������R���ٚ=�+�� �b̠��(3�b�R�Fӽ��N�, E��z.�ZYD��8�k2�^�h���i� `���
�%����:������f�EA��#Z��T��Ĕx��&u+$����0�]T�?s����W�50��QN]F��>e�9�T���4�J2Jq"�x���񭿼Tf1�����5HC�Μ�Ї��e$��
�ikz�k�>E�z��㰞�_��r"
�����|^�0y����Յ���	g��k-'a���"~p�#+�d�� {k=��إk>��l�T�?J��l]�,��3ܫ�?p��	��P�ʸ��Hl�D��L}~<ocTݗ�;ڟ�zl�"WoW=�T+��E#�2H�����]��;_d����>�i��E��u.k����ί�3qC{��,��_T�{��6+^odmO���%�i�EPR��J7s�v�GB��Z�$��"F�ڋ]m�'I�-�oQ�ǈ����Jۧ��������č�BT~zy� ����Ÿn��ak6i��R���P�2��s�������el�C��qZ��4ጝQ�8p�He�M�˂��1{�:q=9�&�dU���/R;�A־�8�����Ȑ˴/���@���Ĭ0�֠^�?�U������ôH�X��6/�2���;b�~�\��R� s'8Mu�7��+�NM�#�^�d�;���"2�����A;��	J���!�p�Z@�l��%�8XO������D3���.w=�@���3�62[��dY���\K��/�>���} �;�][�(�p���OD{�U�6�0��ƙ�4�Ղ!���]�t8qT��4O�YH��N��Ķ��y�H\�{"�v������A�:�?�E�ǂ�f����$�R`����	n%�}�M =��<�d��]���.��4,\��~�%�P ��F�4�U=�@�4D;�[~�عQ�#g�2��<��zG�l����1�t�0�`�9Y�$��V ��W�&v�1��۬��~��������Y�moT]�̶���+�2�.c�u7tu���Cӈ��.qFa3o�ҜN��Ť���'�n���#v��G�����s1(ĭd_$��D�sm�zv����]
���;Qh's֌!�����3��aīW=K�;f�c<��I���e�r�.���ͦ�-��<�E�S�BԮ̘Aّ"��Ѷ��{��c�,�.���|��iV����+m�ޠ�,�!|:����m�	4�G9����"܌!V�B�˙�Ǉ'��%���)k�>���C"o�����"�>���߾���}�i+��8%��lV/��]QRcJ����^�4�)�>�}iUv�*)P��>�[0���( 0�<e�)S[�6�*X�U�UU��$�;����ug]�B�㟯�		��)��)5�oC���2�Z߯^|�iԼ�m�ju.�
��ܐC�E�4��Z&l�M�s���Ag�ҫP��F/0�$��d}�4��ǲ�]%!��I�MG"��D��^�X�\��A?�|���J�p���l2d���Y���\�#t���X��ڍ�Ѕ���ә��WrO��L2#�<���?;�<�w�x�L��F���]*y��d�OL��{�	����u.)Tr4�"��v�#^�HT߿`#�����=�Ș�$���Ő�����$��Q:���/�P��0ci&�e�-+x�Q��(�-�!ǂ��dz(�R8���~�c�G٤�Q����zڑ��a�!�	���R���S7���
���!,eu�0��&�u5��^���-�m����ש�H��@)�E!l�tĠ[��\]x`{u�t�[7|sԷ(��� ��|{fn:�~Ɏ�kR�U��[��й�G9r�b�Fl)�#edU�ߊ{H��K*��2%6�^��n6��M����Bds�A��<����7�5�֑E�T�z6�S�Ve�ӬH��d qw��L-'d{Z�-�L����J3����2���CDǺ��|&�3�u�	P�}�%�v��g+��ޘ�úP�8xh�_���t����f�1M@���17�R�tp������=�����3�{ڂ���tu�PNui�f$Wx�ʉ����^Tm�Gl�q���iY�yp�JL7<P��`�*HD�����/b�'�����c�j�i5����9���]��Y���xTB���>�D8g�\J�6�R�����*� ���$���^�5�� ��n ��_}w�jh"Uz���1��`�:"Y+|����l��,FI���� I��q�j0`��N��uJ�!��Y�V(���U��O3�N�t���୸%V�o�im)]���tD��C�7i������_!����R.\�t,Ō�]aW)�GY��Z���(��F���&W}�O�3��?�w��:i
�C���M��9���A�Y^�=2P��_"B8`剪�ǐ�)V���(!�b����}<��{>í��`%j��9&	Tg�fc/�ʖ��i����괡V���{�_eA�	R��tp�ӧ��"Y���v\
os��<���$s�������?�\��-�)is���S���(ǡP��V3�'�Q����X�<G�����yc�ܣԌn����h\>�F��<-�=�)�Ri=5¦Q$/J�	.=���SO�N;X��HR/�F���T��,<��4��� ͺ7�.s�U�Y���?#'*%���+��]�V_YB�Z�6	��bM��'�v?���R����V1�m`�e�L�m
*23��+-4YHWʴ���G1�X����^���#�� %_)F?鳳`K�
�������Ԯ!<�ea$eK�?��9���'iX��F�S���HR\��A��M���W)�.���L�s�юt�3�#1��5�n�հXDPK<J�i�ܥ�B	U�0w�5����OEI~MVi��S��A����
h�S)����4,r�.�f5�jjldg`�O��ʫ�`,͋�=(�-��?[:�t����Y��WU��DE�9���Y�ӑ��U�r�[��YR	Y3�P�hotR�zԦ���fׂ \��vE���$Ok���HЏ6��sO�/.��I����[#N�\eÞJ�	2̆���Mw@�>�$<��z��C\��������4R�3�#�G��N�Ƴm	���	��2C�#��������A�8�2Р�4Dc ���3�O�C�I[��kUTȗAn�^q�е"�. z�X}}|"��Vw������UǼda��+�� m��`w��MÆR%�'?�9��iI�˴�5���+o��C�� ����s�#N������G�m���E�=����7�LkrҗuO�2#��(��T��g�b����m�'�B$}"���Q�Ƶащ��`:��;D�õ�'K�n����y�r9Y��DIm��S_����>�Ge��df����p1e�5���g3����Z/fԙS��ݺ�����5;�Z@��Q��j@�/�#tZ�S6�eq8�2(0�3੺�v8V���6,�cœ>�9ְ��_�4_��(�U��݋M�⒮f E�[U�Bcj��[�m!��q�I��C0�X'79��y���d���Q�~u:�R��t��}�C�u����W�"1����h�y���P�b�6���ب�6gQ��D���VId��)$6T
�m�6��Ā&f��x�0�G m��P����؉���w�?<�Q)��z��lL8�Jᝧ��)����E��BX��h�3��c��0�T��QYh�_��L�\.2Gu�����m��I��`w+��gW9����]^,ӈ�P�~��mC����v WZ��H@��?��l�׿�� �"��jE���v�ic
�r4�G�N�XڔS�0ř��s�8�B!�r1�BT·T��J��@Y{Dc�~�Y�}o^��Ӂ�l���-�hM�������R��4�Ղ"�S�g��F�����u�!:ҹA���_��Jr؛��d�������U	�۹G
#��փ-Zf|{���ˡY_��|��l����C�<a=�$��s
α��9���OH.��dL��?o��K`��ݷf���n��dִP���0+�4����a�:��"+y2L�F��J;�W��M�]��3ܝ5`��;ݏ{`�Y:9$��E����v*d��+��Z�.�r-���< �O7��0��BHi��9c1őt$5���������Gq2�u�v��K)��}�,@�쮜��$z�Tё�R<�䱷	�迚�S)m3�����ٻ�=9 �6�rh})X�V>�O� �m�x_D�(����������M�[���Hr�x���̐QISc��+�z���Θ�wF�@~)��d�rS�m�Æ����D�du�؃�;��Y�Ȥ�p�lf�\y�8Y����W3�1�@�@�[� &dT��.]�g�A����f�8�(���|�%��y*M_%���ܗ��f?��<�����G�7�F��x�d<�W���2��~{�Á��2/��]����6�g�����ƞ'n�i��Zvj@���}��iq�>�����b�=OWy��"ŜR�x��q�;�M�zrX��|Z,Y8���W�J5K��
�����4��kl��A1Փ�.�I�'�,�!~�=>sҕ{\��ly���D�6�l��Z��ə�o*���]X��(�2F���ʒDZ�@l��:��Rj!"B[}�r�����5�q@ϳ��_(.�r����\<B<�O�g�<��A�̀l*Z���e��3�NYr������U�D�+��OT�fɗ�=GDr��E��d�3�+��3������{.`(#�f*�^RC���
�~U�o�oN�s~�F�+ī�I�s	����%��i�Y)P\5늯�x������j���8a%���Y�>�8�sY�T�Ðw5����{9n��E��#��]D}�UM���$�!ji��L-�Ì�@������Y���a���X	�/�5@��kd�b��%K����oG�,;Bdř�/8%(Ӛ������+@�k�4\
@��Q�c)��Z)6���0b��۳y/�����q�BP�7v���_��A��^M�Vl���I�, ��1Z#�Y�Jp̋��]�i�q}Q {�J��e���{��T'�� �fn���ⲷxf�]�(��4��!���Xy�l�oM���Ug�+�1�6Z
�ko����
�a#5����M�V�dq�r�@XŤV�p�|ٍ��k�$�H�G�U�|#�e�*�DU�yJD��ITȤy��f�I���?�z��m`��`�[n��~�EA��<ěO ���aFޖa��ld��w=J��RpA�H�.E���[�����p�-ޯ_ڣcĬTC��E�O�����d�������:�(�>��y���K@8�P�y�ޔ�J��3��x�N_յ��k}�$���g��{�o%��(��q+P1�N���Oi�Ut�-�u�}�s_;��D�A�?l1c31�L�;�fG�7k��G*���K�:�Ӥ<l�\Sm7u�mXs�7��dص��`ٸ�R�B�X빗ZY�_@N}��]��]ip&����-GN��p�QP���&�(��&�����7�u���,���;���G��!5ƆX��K�[�9NVi:p�������WR�Co����pi�¶jCGf�/pg4%�V5�@��F�\<�=F
����	 �8��D��U����Rd
b{�B���1wJ��s&?1Ll����+xI�w��Y�߸,�	+�3�Ϋ��l��nv���z �#�ÿ�bf���D�6��X��ڶ��1f(g)z@oA����ڒ�@��"ʻC�\�Y�c�~�U��X��z�#��c��&$���i#�9a$�k�p��ye{9Z
�U�'?��`���7�������=!hT��]$jz�����q��'��2k�9�üߗ�_���Y�R�"D���횲����z�ow��oT8��޴ӣ��Z4}^+��}EN�ޓL��ԋbtщ��g.C�u�5��d��I�j�������Y����=R�m[�=Q��a�b�i<�߂�;.����w�ֲ7���m��<((O����a�ǔa��PoiR�<�W����-�TH�.#�Ն�+b���E���3��$ɓ�ݏ��Z	�LN4ق�='v��QZ���Nz�~:;~
���6Z���R�\?b �6���|�#L�c"p&�О�H��r��=	8-��uGI��K�����{��8�Qɳ�#a�RĔ���uE��Lk�-�,!,/� b��P>o���U.|��ST�x��5�C�:��Κ����%U�ŭ]��k��Z]!o��FEt��K<�,;4��[ώ���S�F�t&���J�<��K(�1"TT���}�4�-�X���U��qHE;PSE����b\��yS�5,�-R���꿰/~���Қ˖��:A������_�z��w�"2�gn�^�I�pm�zP�������I�(P�hJ-��`A�NQF�z\����G�7�V�@��gt �0r��b[��ϢګyH"(EU���8Ƶ	8�Q����@��L;��q�\�gF���rFO��\ 2R� 7�q���n6�ډ�Q�nR-��f��N�����) �?�̉Ƴ?�Wu�0�z��+�.�=KVw: ��L��¦�Y\�;��|ŋ,�IQ�����Q��:�k�fD��iY�,�j��?]�����Ų�Fvu�@��a�N��(;�B�V��A�9��)��8��=��^j�9FP��fS��O�����krv�X[C����+��~��� g�n���x���HS�#�F�0���#۝#~_�k.�
�3g��>nP:	����9=U3��rMK�(��u���l0i�<�ΨU�'iEy6W����
�����7��*|<h=lw�U�c�AL�-�6��`#,���*p%�<>�y��,�T�����Q����F�X��b��,�$mBI�ת�� B���_�	6�E�ʒ�{ЊWT��T_�KT� 9?� ✗a6G/܊�yV֟�J"�2B�$3�|�k�Gd�zy"w�O *�餳��R�Rl�m�3�xA�����%`&�wil꣬���Z}.�j����-W�Hw�$��߈�t�..���s�*�p�n�2�{��`�Z��?(�gP�F�&S�{PKZTj���ۤ�Q���>(T���EǏ\h��瓜e�5�25ywJ|������K2����]g���q��8�4��x~g6Ɣh��c��B�ũ�|LX�Zc�-"�;M�D�#���QgʘכHN�����5(hċ�ԣ.�f=�6g�
#;:ا5�W��f��j�-^R�e�y����Z�M��Ř���|4؇J��
�+�}��}���p��ڃ�0Ѵo�H��kp�����@��� �"�ۧ��	h'�E������å�#UrV����
�qI����H5��.|�\���=��ĝ4N�{}.�e�31���e !����m��٤���8���N/
Mw�'��i$�PO��RJ�O�C{���]�=�_�eq���hH­�O�̈��ٴ�Vz&Q���ڦ�Eݟ�G�P܉5\�)9��6?؞K{u\0f�"�m~�Y�A哚R�/Y[�O���H�i��6p��M|�w3%�X`0�3���#93h���8?���t���=��6{�r��e���Wz��F|��� �SPh���E�4S2[�ڣ���TG�S�)p�g
�ϛ	��i��N"�W7��;��$R�=�jEX
jmHO�K��D����1
䍤rFm\3����,�N�S�1����`�h i�i'���V�GeO�����{��Y=��:�0A#w
���J����w��� @�$�F����?� �O��lƢ>�˯�x9B���_�Lx����9&�^�5�����;|~�>@1T[���v�%�M�(��c߈��0D �44���'��������{�������};-�i���s�4%&��r��L�B����Y��ܲ=�|Ù������R�����B��S�v��y��xXm@�����K��R}�+P��zg���K��{C"����RO�Lو��/_�;��5���:�u�����a�އ��e'�LT���o �c�Ӈ�y	g�[(��c|e�S
u�i��<������������<� �h��2�x%)�_����b|��}\�M��)� ]�g��1V��������KIY�jTuμ6�����;�R���Yl���[r:)��Q@w��T7(��x"Lm� RX Q���v6�n�Vߖ힅L���D�Y	��)?����B�%��h(��cj~��<\b���h_�S�>-��c�����O,��G�H<��{��d�X�! �;@H��I�x/�4�d&K�`�Vd{]y��O�]��=X�#�Lz� ��/�:>�f�[���q�M�����Ԥ��bo
˘��x�.�&�^+ꤺ��ۓS\1�؏�,��T�zn9��;4~�U�5SC�0\�E���������jM��#W�×�m��Y�vRD�Թ���V��ץ�p���d�$)ǆ�F����eoظ	3���s$��n����@㱕��x�+��΀B�G������]!�Y6mYm�|NWn��V���f�@�1L��=�hE:0"������T�נxOV�%%l��^���&���"�ߠ�Lk�u��뮥�^<<�+��m�����[?..G�(����Έ)w�3%�]���T��㿬��gM�<hF��6�ġp���m��i�o\ty���Β$P��A�	b��t���7��WBx��B���R&Q5[����W�����xoa�e��Վ�R�������� �L��T-�L�)?��aXw��iG��7���}��ePu\�i�X��Սk��PW�����L�u�0�>��ӓ�Px��J
ʛLHF�<�K''�F��sK)��h��ғ�dr}���u�>I��P-p&�Z#��U� ↹�m�q�CNg��J�.�)���R��57:�K��P�1x_��N�`��k��~CL*�C+��m�u[��}�s�&�FS� ��+��2���I����t�Q?���Vq�/����T	�-��.mT̔O����n��A�[��b���Я�c�-��I�t���s}��Q�fm��zV:ۼ
- �	"��g��[4����]��3���
xx�S����_H�J{M��[�������������(A�1��4�C��5���|�5��E�7ɳ~f)�	��������{@2��O�2�~��Cn��d{f�݉�PP&�&QV�4�Pw5���xx��|wE7n��z,�R�q�7�n"�1kW:���	�]�;���=�+24u,���[����י���o@,"#��Q���7�!����c�
zG��?�p�q����t �«ǔ(�ck�/-��BLQ�ed$S=5,��=*F!���3���A�c���� J�u���AѰ?L�J~S,tW���)�a�/�CrW���RRш��{�H� �J��ķGE<����V�?{k9�)�r
:.��m�]4?֕r�M������ˬ�c;�w�uw||�K����#�Hpm�b<�G_��?#�=�7 af�����@s��cc�G�����ޙG�@�[�y��k�b6�;�i��𼝮G�i@O�������*o��,���0#*���q�h�v1}��#9͝OٯϮz�AedE�N�Z,����k(z��֐ܴ�u�૦�����`׭��i��)�΢
k�r��4B}bo�_��Q������0[���t×�R�U������ƍ�����J����s�k����֊�F�%	�x���@ԩ��<Z.~��ޜ��(�é�� �%l�X��}�-W}�\�f�t��_]�pV�.�+��n���|�Q��"�v�HS?=9t�ke���|��,.�J���f����V�BT�T�1�;�wk]����	��bC������kdٕ�L�4����FH�^��c1�憁��+��Җ?����
������n8hD��M#��7�vF��� -��R�꿱H�4��Fh���'Ȭ�׻��.�����$w�hv�}�.92��q�2����0�P{kz��a�>]�OG^�nC�f�qo��o>���M��~5`�p�A��gȥ��%���&-W���c*]q�>?;Vzk��B�_:�q��O�&k�V�ҒgeR�t؝�(����}Ҟ��������_/L?���&��p������:�ܟE�[�?�S���Ug8����(`�3���<�3�D�M��v{U��}c9�Z�*C�[T$sz~�.nz�XcD��0���v�ԬƤ�]�5��w�k>���s�a��ق½%���A�ga,��q�Φ��áx��Y�oM39���(��6��RS�Z�|��ad��9ȼ�r��Ȇ�ں��u�kMwl���V��ɫ,�7J|q���
��K�Y�O,�'��7{�R�**-b��RE*��b�e#���p�0��3 s�Ӛ��r�����G�3�l@��AKF�{��`�ң�Ι"_��`}����.��\�ɠƭ
�Savou���m.q#J%7�|\�|'!nDk�lŭ���>[�w�ţi��O���B���q�$�tEL Q/v�	��h.uDC,C�	�{r�Lʐ�]˛��z��&5���U���2k�Ct��,M��7h���tPMΐ���)M��+B���,P
`n��`
6��u���5���5�J���$��UzH��<�{�% ��G��"�8'��lӜ��	T�0%��x�^6�xo��A�XH�K)����]�8����c͒_���D�(O�/�2���C���3��!wS��k�ف� �M�kQ��g0�4���7u��o:�aPAltOkz�4z��S�ڹ�l�h<r�!���\�n�lV`JF��TUrg���n�}<E���%C���3�b�����Rx�e���8W.����r�K��v�����/*�`�K;�ZACm�%�@�DR�M�#��g�~�Jq�"�P���`�MX�pґ񾐂g���3�l6����J��}���:���To��j��8�����ee!XW?9N̠���2o�?ᬷiE��y|G�~���K��kHm*�9A��?>IǦ�ՙW���F��������!�1j���/pn�,⦖�
���J��a'T>.!��/���m���c�����̡���mf���.I�E�G�M�xa8��=�+יr��S����(/0�uvo�q��7͔� ��i.�M�[�]�؋B�����u��.�6���ǙE�2��h: Kq��7bB���3���+0WKi6rg�/R0#��ϺQ�oN�J����fZ�?�'Rx7K�O�NR�'����]SV �YԞR��8�@%�D#���ơO1�ܥ^�nѴĈC>i��<��:k�e ��Ϡ43�]~�.�D:P)u]�/)�q��D�v4���ت/������ey��ʩ���&�O9n�@�� 6F�&�$|�uバ������L�yu?S������	��%�B���>Ⱥ�)е �=h��?#5�o�%�����v���W�=�h
�j'P�?�(W��3칵H�B֊0Ȏ-+�I�����re��P�{E?�%�q��ӣ�_I�]֧ljt���@B�@<^�b6hD�E<�9��4����:�W�h��~�ԑ���B�{۪�{-_��_����L��q�3�T��h/�we<����fnu�~�J.�9C��#ӕ��#+̣��	e$8C|����O�֞����l��h����i�	�y��Yi���etlL��Vn��J������*�����TY���r���:��Ø\����i���FI`��\	���\�t�M�5;��y׀^�%|�[lP`�����6���`�.u�7^W�(�y��7�A�G��>��ӟ3%j�K��U)���W��rE:C�����u+�6�V.:��醈����YLz�ň�N���h��o���3����1a�����>C[�W������V�)����UT����hΪMy�ͧ�����f�P��g�K�)1r���C�`	���[�����;$��,%��x�@��,An�q�4t����o���>L�� ���RU��"�=ħc�0�F%��{/m��p�ag;�W}.�9�|��t"���K���NsG��TY���|�\{F�X]��k] r7�E��Ѻ�U�ƹ���;3 ��U��Wz�f�,�ÐBe����%���ͽ��,YNS�	�����OVvp(L�[k����HeiIg8fՈ�~���7o�}�/=Қ+ꏣ����
2異�6�MJ����6�0�Sh�ǭ{�sǸ����3õ��&�xSg	�a:��Yo�	+c1n/"S��h��%�xׄ�\�Ic�Q%1%y�-"�!���Ҩ�F�(��k��U]�3��p�6 c����](��CZ�Sh������Gi��C�$�j5�> w����/̉(li߈���o]�OpmH("� ���3�/o.�#�YW�M��ץL;i�� �2���f��g���b'�j��+����n0'�߸X�N�S;~e�QQ����7�x�e��}�x*s��S*u*����(�hy�v��[sO�ta����κ5��r�*fYKrv��x�aJ��5�M��7��#{��qC���5D�x҉�����ox�C�)�L�>��i�:p�o��0\�4��ch�2
S� -f�v������m�:�,L�T7�l�~qB�N�"��D��23���-���`�C�z�t�ݕ�)��W83���2ե���[r)�n�e�sӆr�c����AήL���v���Q�!i���I�&r���qԚ�#�Æ� �ĝX o�-�ڋ�����`e�y��3y���5Y����,���2C,��j�I���d�Dz����yi�w�)��Bw��x&�}�.��e��(��M	b8��?�
�����}^�[�f.{O�#������Ã��:��؟bL��^�(M��Eq��Ȣ'w�{��*�?�;�B���w���-5�͸d�����·���iwQqE��2�ˠlh�S*�-E�7����R�����b2�m�"ӎx3��W(�'�t�����0q���er�Q�XR������@b���\�Hp�Fi�0Ƿu(�� OI B�8f�U�;/���w9R$��"�.����`��I/�A�8;����D��Ag�#�a^ɼg�����0����;�-��kACq|�_^�G��+2О���{,���Z�hz<�jWIq#��霳YJ�ʺMAW>�Mh��{��#�:0�JjR�9z����©j-Fb$@3�K�J66�����쟻�E�|x��nR�):��W��U98c��\��'k���	/o�D�?�|���?�i�sQ��P��wb�5���ΏOő����n�[v����6^~j#��j.L�<ШOR٫"�G\x�H��oˋ9��|:4��U�� wFS�227S�n��!����j$�L!ȯ��B�����N�����.�����W�����u��]�p��9e/L�\���Vq7�����[�k��%W5��k�xy/�������d��$"���k�H��+F�t�[��c�If$��E��<���F�h��?��s.ʺ%4��'&e6=>#�B���-�}���'�
�^��]w)����3JS߈�{�b���W�� j��,��}WEg����݄:�.`�@8��f�i�oM�Ϧ�Gw���F;��a�O�E��>e�L��v���fs$ l6^���Նt��*sd:�\Qnꓬ�@�Ȑf�#�`��vABZ���k���0�%?��߽�S	4l9[�9u� Ζ�3I��]]T�} �]�m#F�nN֫jK�ѽ��t"P���@�:�;�� �P�LN���Ͻ[��E��Җ�w�Z=�����!]@�8���w [�>��b�1�@��D,܇�=
um.�ri����J H�_T7�����r�m��g�!��r����/&��B�[�"����Y���Z���Q5$�=��0o-�x�|�t��:�����Y��q`beu�Rk�*g�On��7�xvTS
R�x9��y3s�\F8�{$ҰZl��R�V�tM/bSsJ�����I��l%�5��]@¯�`��&F�	
%���+p�y�#�&ˢ�%bf���s�4pP|��?ȳx�)������ǧ�ޜ-u�ٺ���n(j�\~[>{v�n���>^��R��&�<�N(`����'�r�}DJ5�<��;p��D�S��
(	p��$�$�0���ۢ��*�9L\61a�29�q���M��ݟ��0��Y����>i��;�As��>Qj�1�VT�TP�����T���?�f.rZ6�ѝ����4A6���p�$~ˢ̫��uKՍ7EV�lmP��ڿ�c|H)k_ ;s�Wje*|4��R�Zy`|�(F���9Tf+$/)��3�m�Z���(�M�*{�uG�Ď�uX�5ψ�c^S�0�$� G�5r�T)�Ώef��%�?���0O^��xS`�.-�]�wݑQ:P}�+��x��78�W�ʢt��
��r������U��*��9������J��`�����v��3T�5�I���n��)���2��L�wTp.��[�m���$��qK��7^e>Y�%�%��b�Kl4`���ٹX0AH,����Σ[��p�6:׳X�!%K�4�$���
z��P������H��:M�vxg�K 6�ڛ�Y����Ǔp}<=����Ɲ�֘�lޖ���>c��`_b�lY���T��-�:Y*+QP�	��s*�X��9<Jb���һ�H�7> 8�sǖ0���Q��4e�Q�Lh�v��>[�:�M#�R�雑zAq@�]�7 ܆u��E�w�LW��Tųe�2��^"F��;�d�S�|��s+�,]�nyp��l�Y�:�l�%#�EWR���A����vUU�Y�L������=�DۘoTr����Y�0���H��Jt�V�ќ������)ů.q��r�"�O��,� �ֹ�����³-	8��d<I9� ;�Gi̽�M6M:1"ڣ~I*�
׹C�7Й�Δr�'M�I�S(_
�B�OE����}���	���}(��fX�gr�v#/FIg��PI�������ȵ9�gd��ھ��Ts24�\��ū7��+m�4��f>�P�j��qMSn��`�$|�zp��Q.I��b�M8oo1��ܶ2��7��,�S�L^%'��WZj��]��-��>E���]�w�V��[��TX[���O�{38�U^����0�\mN/�"���.�}���r�I
�m��D����)�2�k��Ҩ*�y�(9aO�ǙB+x��b�wƹ`wm���!ۤr��)F\����C��"�$���ٟG�&���<Z�z��t�;W,�)j�7&�+�Vb�`��|5x�4�Q���r�C*͇�A�ۣ�[���Wm��Q�'����Sp�����x6n�cU[���jd^7_4<tE�]�!�P�n�n��Fb�$9�}�<��- u^OF.$�N�i�B] �'j%��8�J|������7�4T-k��L��,�3��h�ﲈ���7�������~5Z��;�u�E����@�X��p��!M�H`�Z�7��'i=Uu<�0�U:E��"u�����[�����,�a�UiGGߪ�ţ�*S�c�,>�iR��r~Apۓ�����zCΙq�@�ŘQ�ц�zb�q�� ǩ��Ol������w���}�E	M��M�B�nQU,z�k�g�����C/զ�sI�S4��{��U+��/���N��>�ȣ��Ũj�����(?��V���g72�m�tc�4=jD���å托���L�6�_�Z�p�I>#n��j�s3C�&���84���,Q ��;�T��gToGhU˹hH����E�B��u���k��)��03�{Ӡ�Cyix�C�.�v`���x�ж�[�Ջ�]cr���ˋx�<�J�E�+D��7�!�q-[�Y�k܈�l#k�#W���x��L���a�Fp�24{�{�'ı�T7�"���>a�In�j�}��}���
��(��6�Z��wCU�B�L�YD)�\���[�#*-�Gy��ϊ|Ƙ����=��2Ix�d�:vaH�@m"���{�x��nZ�S�YΒ�����.-�q�i���w�jU<c��n�r�-�Q�NRe�p�AD������rJ�g=9jio����7eR�1���4�#Ũ�I\:J4x6k��CS��06a2��j=D�Ӥ�޶�Xr�NV����M(�=2xWGG��އ65F�B�8�iF�����N6��n��|k=@��ۻ5�zN��5-f̜�.*/d z0"�*7I$aIu��W+Cr�_�ٸ�2|�nR���΢|���;��߇؂O���L�#V�?(/";88���K�%u������j�9�_�z��e H*����5��0��2�)%v<%��kUD�Ն~�t�7��ڕ���NX/o��'|gߴaxˎ�)�H�K`B�|�n�-���(�T~�&����9f6
%����<�&rd�Əe���_V���C���}�@s�w��2�&�B�A�o��������,vY�4���^R�	L�Ѵ�?�r
"@3�&��'%h%@}��W�D����ca��T�b0&�D�P��>Aȴe����4�|��R�9){��)��'��V7�r?z�L���G0�`90G ̱���w8�v���JD��h�N���~���#��&m�Z��)�e ������+3����Dg9���%jO��=!�;�y���&�_������E��T���~J�Os|���P����d:>�4n��|���g��ӥ<�'D�j6��n��S@K5}�j��h�α`}	+6��W#嫠�v��{�pޟ��Hbpz�I��k���K�I��̪P-�$$�CA��Rz����y|CҚ��话�.���?��@a۞��4�n��Ȏ~�.M�X8%$n Oyj�֛�&��9��1�\��wu���:dG��\'�K~��Vѥ/�g��&>Xnk,v��8�|��VlN]qڣ���$dQ4���0Zz�k�f�Ԑ�s�L2	�xRx,��Q�z�/^,�pI4{s(��7�84R�T��R��5/'82e�"0�Zs���nm��޶���1���V��7�ť�"���A�!���;�&��m%#��EN��nZ?	�0���|^���ҡM��.�f,��� 0+1�sX���8��j�6O�.B 6�˧�@x��F�X�00��X1�d�Vާ�W�7��@������ݣb]���I�+?�i�DOd����a;��TQ9�F�
��Ǔm;=)�(� ��/6��G+�Xۑ1�U�'~�&6�
v���ao������o�c���1�R�=F�/U��{�u(e.�|'�N,2�q趬��.v�)/�ߘ#�鷣y"}��^�I��D����-�\��o��C���-��zPqAT��D[Q����Iol��z~پ	�$]����
/>Y��0Ə�|m�\A�H%\O?O�Y.eŁU�>���斏�е��N������<;��%�Y�AD�:M�K���p�&P����D n-�2<�i�Ḱ�У�qLB�{��
_n�����?�+7�u <�S~�c�m*�.͗��ϧY���z9�BK�
��"�\�/Kn���<�@NFY���޴��=C�F�3��?XE��$�	���#DƁG&��S�σ��M����s�tQ���a���E�	���t���f�F*A�;�2���<�GF❍jR;�{���B�R��BԚVQ�\]d[�pu��Uk�}����Z�X�U_�����bȩbl��0Ǧ<�Ѥ�{�( ˴��_E�e��Y߾,��żM����� �$p�]�)�k����,�\fdI���	���lB�X@}t�9r@�P��Z�f%0��3�M�8�b�\Y��)V�� g_$��?��%���F�4s��0��D9f���B���h�Q�Y����s���0+k����P��z�-��es���L���}���
�Q&�,�XN�-�:4�����oJcVlz�)�P;��45ӌ�g��	GN%N�I����GRN��������=T��M0�f��/��������?����-}^s�
6
O��ՂbV}37�{C�V�b�f�(EM	�����h�{�yt���ɨ.�%�Q���X�Z���xIC�e�g�Il4C��K����bf�R�*z!<'��Y��_J,	�t*qi�����¸Q��8�a�	~S���>��3�cS�t��<h���,�;�M���K�"�/�+�)�6��<�^l�e�s"�H����G��m���s�Sk|F����FE �M��`(e�� ���WE�^�^*�'!�AĔ�X|��m@�r���t�3�~܅�޵������
�C- �d��0�E���G��<�HX�7���^�ڂr�v��������c����h��Nչ��|�?�c�xG�}��ľs�Dt>Hh�t�-��ߍ#�5H��-S-�.( �T�Q�E��ePT,�1��8'��ѧE�f�є�H7�k��P�f �t7^��披8O�.��%ߧ� �Zb�P��`��9�k��K�( &.���Bb��j�������Yx�b�K��\�G�M�EN����A �@ �sF� ro��<3w@ن��+}\�8P��o�Z7���<��m�`0�����b��/y9�OX��_������
������yk���&�4;n�M~�p엾^ٶgE���z�ׇ�J��7��U-��QY�.��|���D��l�@h�P��6nƩ]��36Ж��k���2��a�_���)Ip�QC��ߴ�c���,�v���.l�h�h��^S=Lx�}�'� 8-�d���e���;Ttnđ�G�����z�'g^r�>������<�;J&��R& �����XL�1DWJg(��EP&��������w�J7�r�򕆗��ٔ�Jp��Փ�U�H]�Z��u0�5}זi��^��@���դK
�C����&�^Um�i?1�5���Y�]�_o�#�ex�$�X�$�a��[����ݝ	f@��gÎ�
zJ�q{׬��@�4A[)�e�%�FLh�A)K���|���g��$�CX�.~@�T�c�Ũɯ{����J'_zm�� I�<�����Zw����w�3uY�f�*�@������_ٙV�"U�Hn�>�EhRgGKd� 2w��|
~��V9�E�����w#R���I����e$;|�n�~��\ֽ���|�g#I�����l�T5�f#.Ȇ����Ly����4<-@d�������tՃ�͚֟��-H�k�;�����e�a#��(;&b�E�j�s�8]�o��a�m�e�5��RS�'%R��8l��3�Au���1���{��މ�t.5���w�� ��!��C\�<?>�B�x>u�L�MDR�����H�9�a��pR/�~���
��H�<�⌏�8�{��[�"��O��!��
�vY`�o����X��J֪#/��\&xw`z%�b��Km��U�%:L=[�w�:�����|���9���b��8����9���Y3��	R��]����[��4y����E'*��x��'}����	Bm��Z���]������{�G����C��������@��M(������-w&I�	y���9[����`]v�hRZ�F��̪�!	^U�`%�O�OsŴ_���}s�A��i]JY�z�mvi��zb+�%���:�還�c1��?���LO�Z#��sn�������:�3��?jo8�w�p�^���a?�p�cuk�w e}��fq���Al�%����\�]�W3��q��I�5�;i�-��H;�L�\l)f% !�h�x�>�4� 1I�§2�3)�>�ባ�a�&7��^�Ռ��ZQ+,��&���]���n\"��ML�ּ��Ο~�Te�����u�
�Skv��c���a�:�7�
�l���N�F�����0w_l(���	�v�C��T�V%��F��4&�ϋ���ؾ�bUM�1?�aT|��E���)r�o��j��t�6�K3d`��������p(����e7���;�>���(�?��j�����zd�_��i�=�C���� E�/�jq�w?��o|w����6���aQ���I�����}���]��x���F����G���A�Eu��y`]G��r���Ѷ��J@q�p?�E��s�v���D�}����ֵ�{w�VG����ǣ� y�\p���ĝ́����mt���_�LW�M2���ْ i��~����^���FDL"HCY1x v�OhJC̢��e��;m������ѐ��"�b`7{[�=�<��X����a��%-,��>�m�W�՘@i��m���5�$���i؆m@'L)���
rİϮnertv=�mk���f�.�U�$@�ITQ�G�GNO���xk�v�O��Q�*��h� ��=�h���|�x��\�Q�|c�B�pK���ͩ%;��
P����V�1�"^D���+8�R��vt��]5�`��=C^:"I;붔l�I��K�Lh���D\�歧��|�ٺG�*���@հ��<8�4|�C(i�{����Z��`�o��S���\z$2��b�՗���-�~�-(8�9t(�Z�A�Fx��_d�\{{,��n���D
���="C���\f���zl� �גyNN���4Fs�g�̉�ͤ�"o���`*�h[�qWcA-(�������c