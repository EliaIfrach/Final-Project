��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
~����KU]�R�X��2�T�V�t��[T�v_:�4��q�Ig�>���[bD�����^���s����ݑ$��7��1B̈́M���wM|-�TeV�( id��k��cXP�Co�3�����|k��$���a�:;�97�{�K�"���Uk�	�) ���6�K���W�Z��u[�K�t�z]����LȮ�x��WPC򟂪�վo-�OS��º��kjS���@Ψq<n��i�Z�S�雋�f��Z�]Yz����և�c�{��?4�A��NZ�.��y��ʞֻ(�n,�e�����P*�JP��}�^|����E��*m!��eR�����{����)�F�GLqd�-�u�) ��Y�U���?�3�_	�=���yz�P'�����闤=yfߐ���	�P����O���N��Й!�u$�kN6�I���
!o�#��K�l���Z��Z��?ٹ.�j��h��3�5U�Xg�>c8�KM)���}��Vٜ,ǜq)e��_�w����8MVz�X� E��JY�"����	��B'���Q9�ͯ\u��@��A"������1/=����~$���ۘ�8-��1|�Æ�`�wzܟ���}O��� ���� �k��� �x�_�*�0�U�#D��]����h�@��qd!�~���X`����^����s���O:3T2�kk�C���O�ѕ"[�'!��yF�}�L
�%K}���P-�'�!�7����O��#�I_S�׺2�bDD+>64y(Bĵ���V ���m����u��Zw���I�2.�iLw�ݪm��}����Ր�Uܩ����W�(F4�F���N�<��0q�38�3)�,r90g�m�w�Oݔ[�h׋�X�q���]���b�c��� [DEV�,$=�%S@�k�f#y�����-8EV��/Ν�}C�t�L��ol3�CA<s:���� *l���-�yOj��1�sJ�Z��t�q�-��=l���p�_�>_����oRL)K�^��q^���r����]u[F�W��ߏ��v���y�R����|�`h�j�d�\�1-vC�r�Y_�>ɖ�� �7c���z/����ޡ�ݝ�rP�c��Z�M�j��`\��,&7y�:旖I��2���R�%xe�{�.�4�
�4<3P�A8rm����(-��F�	O�����E �_��;�R��:��܋pA���.֨:��O�ҁ	P�I� ���E�*S�_��s���p�qR�y��-��=piU1�l�%x���\�M�>�L꾀���&� Ob㔃Ulf�A��1�G<	4�y�cЌz(Z�@{/�9���#\�Sh�%砄�0	���l��
rW�u��~��z!'���_o�kZS��ܔ�=B��_�Ѣ �럢$Mf�|�{;�o�F��C,m3����$����2��	A&K�3y�����V�'D��PEn�a��}�F͎��R1�V&�-XUYa� ���0պ3�˟Z��j��
���t0�)���Yaڣ Qi��b|C2�V7�p���f��x	��T�){>L��5ȫp*�?�ǹV�]<D�K��i��X����Ƙ(@�_]��l>*�5�k���aϘ��R	��Ž�
"2ȣ��MӾ�L��[~h\!?��%3�'p�i��P��Y�q;�ѩ�X�� |:�U/\o��)O��W;��^��D.^p������u���F�p�69��q�p�ß�+Is��V�WD��i���1<#:W�e�a9����dZ�VR�l T�9~�[����_I�+Q���
�/�ه=?��m-f��ȃ�w�81�3���M������V(c�>\Q�+�� p�{�y���1O���\�m$I��R־��W�at����L�z���Z�c��F~��DyL��[�7����0���B����� �6�s�LS9�`�z6�Y2g��a��	Sl!����m�Ӿ�G�%޲3�(wy��5 k�}�	�$	�Ch�GQ�B�8���n�T�5������Qc���"�تR?����g��O�0.U����,��91��~�/��"01�M{��W�s�ss�c_u���j���Ʌ�ʋ):(� T���ڦ�&���C��o|}����ԟK�SW�徤��?�
/w���zU��)�H
'��7���7����m��c��� w�ƙ2)s�}{!�����K3ήh��V�9��nh�D�"L���K�<�6X��G�>%v��$�pB0эTh��*{��d�a�Rq�BM��Ǔ�J���;%�4���t�[*�1h�_��B�h�IgKcAٞ��L;���wܨў�S��:X�s��B�X�w/B�c���V-P!�d}�^51�2F�]O��.wy�v>��(o�B<.��j�W?Aw�zg�Ltbfq�.4C�	p㓏�q��nN��x�l�orң�Gɂ� ��4'Ѱ������8+�cmĢ�e�k ��,�3����v~@Jڲ��S�.UH����n��5)'T�ģ���3y�����W:1��S
ucV�tW2P���r��F�]����,o�ɻ�m�(�hr���Q������l��V�⠀��%m������l����r(���"�)���l\I��<Jx�>�V���W��C仧��}xEeq�� ѷ�д~!ZL3Re������n�]ᖎ�m�D(�5�Th�A�A �����U����cɿܼA$�{���e��/ep�Q�#����%B�n�3�H��Kqe�f��Y������v�A�{Vm��jT����wr� ��	��&�~[X����;j�b��c�l�Yא��7�{�ug�O6f�:)2����ڦ���m2�n>CSK�K~��ʫ�7J�y� �7r��ݡZ�jMw�]Ĥ�t�Ϝo{�%c�E9�~p�#��n:��_=)݀|Z����\U��L�-�V:�啘4�`y���t׹��T���FB�O�7{]OG�w�¯�(���E?�ۅc��M�k!n6���	�L�ڿ={�:t��s�N��5N��^�z����<��3хw���W�d��v��
-xZ��&4+R��"!����E��i$pDV�㿤��^�׷��F#gp�Xmv3m��DѤ7�|5��X�����l����JFcv���oWUtq���{o�&F�q����{L(�z�>㸳���$�B5ɶvXuC7�rw��魎?��wV�(�0]J��+1�;���F"XN�*�҉<�B�Q��34�p��w��*�Z��p��u�]�Z:Hފ�N�T���.s_��Y��x-���"�"=��m߾���B�GiAL�G���h�~WC�](��{^AM��G`�T�J��h���6���}�%N��I�����^�R��*��֔�C\U�s�9�������(��,	N<u�~s[t���Ѵn�iF�6���eEO\�rt[�f���=\6�LH����@�y\����N�ֵȤ�d�����Ŗ�5��N��H|�%s��Xm���:6+y|�8��k-�P�Ѹ���F�N�r_�w�7�����=�����|} o�	T�0�)|KP)��OL��ٿD��#~C��n��A]b���W��g8c�