��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
�������>g�2���ۆ��6In$�[��,)E���������R���[�g>�6\�!L���G�<�z���rݲKG�L�p�3�v`�g2og�3cп���m� ��������{Bṗ�6�Ʋ���LQ�T���U�Z4��(�Ϡ�<x�>j���^10arrh��Ɂ9�wKũ�(Qul,7	�}s��6��z/��Y�Ҭ�b�ԡ���1��ߌJn�8����E�	h׌�K�!��	vXU"���:��$Y��T
pl,��N���bJ������5��<�i�qM�Y�����e6�ҍy�m!%�2&�	�#"C�S�_� qI�Oh-5�"�ّ��w����)e��O�6g-��W���w��7�弣�mM�Sx8RFW9��+u��')I,_�.���Bd�a+�����J=��	u�kG0Xrm��6�Ϧ���Z�9xK�<���MUg�������
�~�Q��Q�A x���X]�����h�;ѝ������IU��6����bJ���?�����\)��D���m?Ǔh�ĳ�qy��[��"�*������c���O�8WWBՍh��p(�����ʸі�9_����m��,Ӂgo_r��?8x����u��Z�ܦ�pE&J��Q��G���?��\�t(�� oR�
h)s�OU�6p�������g���fe�C��u*޽u^Y*0 ���G4`��bL �U�~��4���Ts�T!Ҧǰ>��_Ci�zdh����m67��f��wv!>������o��0��b.v�=��4;�G?Ut�^�r�!o�e� �D�\@Qޱq�'c���W� ���/�3?�>�;��ѷC������0=���ә�m~�¾�����9y�<ZЩS�,���*v�\eQ�GV�����rfr-~��BuWQ��Y���s��>r����5��쀬���x�髾� C��nR��W�s�D�^��of��� �����܆�	�ܭG��p� H�骉��������@N<ј�Z�B��d��/��6�B����o<�sGa����\�,L��o�Y�h�{	�Ƒk#�s������hb+�⛋_�*����8'Kc�s�Tf�0]U��Ǘ��xhS$݂�*����2��%��8��IU�+=���{|`HL��.�͕��M�sE5=m@��BN�wj�/�u�nG�E`!
D��3�E/.<�T���h���M%(��8F� qy�� f\?��h�-t^޺΁mܡ��2�Y;6���J��+�``��g���`�{��EN�}�Vo|�[/қ
g�!x/-?uLG|چ���Wۣ8ȹ]:�+�ct�������W��i{8$ �����^
2C��P��,��#���.i�����rʡ깉�c��T|�;�7(oN�`�5 ����p����8�wEB��u{��O�h��'R"�&U�+�m>?�6��P�#���2l"��;vt��	����v, ��k��b�y���q�ݢ�Ms26"��qEx�r�ۗ�di�p�H��jk����G]QZ��&��<��Qq*޼��8U
�E�n���ؐAg
��D�
+��.c��4����3�T�ϳ0 s��.���w��m �\�}[T���o#t�8�9{�C����b��sW�n��<���
��j�jzo��ʗ���7��&�;���鑤�aݮzQdeD����LV�q���I��������7n�!�%�
~���&�<Ѯf��-�@��c���,)�h66�Km�����<���~��eϔ�_�}��vĤ:/_�3 �y_1��� ?�*ރ�\�{��э9h�XW�,��H{FV���U���e�T�����~ܐ- ��`[����g��+-(��)��Z@<DRC����8��V,�쇍&,��;[���ݷ�����vO�I�=y>��\Sև��;��!!�����2W?xEY-���^���gɣ��ڣ�e�p�{�8�����a���i��-�-Z���OB����h���ƊH�^%[�zޗ��c�3n�{���v:�T�Dc_���Ҳ�@=������2�	��r�Meg�������.�\��1Q��B�}�CN���n���&݊���JH	g�?���m�)������8|�$ޞK��gA�%�wȑ�����#Jw"�]�0�4ԉ�*L>��<;I�z<y�s����k���$��sܽa"(�_��DP��@�w?� /�W�S�jCd�g�W�2�,�1���PO����J���{!:P��MMXA���@�o^�O.��6m6���~�F�Ru|u�S��̣���K���<o��9�QYr[㌰NK��n�z�V�-=����ȸ�
$5��9��ia�ҁ��a�@�E��2����@򠄏nJ����5��"���5�p�3+�rc��ro�9�
hV���^J�)k�[���B��d�aK�j�7�;�lFHʒ�����o�T�1�E<������<-, �O'�b�
���4��?F`�Z�6�w_B�;D_�J�|^Jp�t6!Z�vxr�mqO�C4�5g��ԍr����r�?
�����>$�6-�2������J���F���9��a�W����͙��R��6����#%���i�=�����-C��g��g��v��$ĳ�}��8�a��9_c�X���5�yܴ\#&�u�&ΨT��L]��xNstF�����3sAgx�i���.�4κ
����:D�3�]h2�j��+z�2y��g+P��yQ��%��Ka�9���I�rD�50`�N��;������?�:�\�ˏz���f~Їj	"H�Q�qQK�~SN���Y$�c-	��槯��Kg��6��4��"����@M��"(�.1N��Wr{�}�Fr�E039P��_l/�2�h{���V|DgH�u���_��JVT�!�O�ǟ�{ZhH�h��m�
�7l`�Gi�(�h�2Yp5���N1Y�&�]���uZv����\�q��|I���d{8�
�8�L&�n|�7p�D���'��7?���MS`�"�n��K��U��A�?�*���)� V�?���a���y E�6+��l"�,:�f�|[�K��(��.h�k��7i&���|���|�-8`�n�����!W�w�v$;de���G�%b0�6�\ ���6G۳�k0���޲�j̦ƅU��	DRP(Ϙ��I�^&2��}m(
��Pp1�:Ť3����-��$[�͹��E�>��s�X��k�=ȍ������`d�3\�z��\��Kp�xZ�b�m��_;�^�/#4N��r-��rpR��j���I9!)���ئ�-I��;T,\
�-,��	��C�:O 0����eV���ǡ�OU�v�A���Yi�Q�fA?|-�����᲌�U7�{�Oz!G�q��)�����;����P��z)� (*:"���C�a��������?���aσ�-�Y���@!aG��J+�(�ͯ��"�$s�s.[]�������QB��#O��l(�K�ǔ$R�M\��Bp�]�~T�iӃ���a�I0�y"�@���0y�[��H0���*X��l~��Z^F*�5Y��uv��[���a�2RLޏ��b�1�t�����Nu/ﾞ�(L�n����D�r�p�aOBٍ9�w4�hI��-����I,	���-r@��ݡ��y6�Y���c����A��WPKҴ����N T�l�X�ζ��&oe�W�x����J��*,4+� ��5������ٳ5>�Bƾ��:��3Ň����G�xix/�K�ˢ�®�����
��z�LԺ�������=�lҒ��An���6
׍�^6s?�΁>
����������[��ܢtL�C4ޔ���Rz'ʟ���OL��r�D@RbN͵����h�O`J��K�Ό��a�ښ0q�=.e[��rǭɏ8�~������]��^S�h=\���0Л�c�(��Y������|��l��m���]FƼ��k�R$��Ne���7=P����V6�\�H8o�V�i�s�`�ì���~@@����ubߧN��y���d����N|���A�C�2&̀:fnhJ�K�#<nX(����Y`H���_���V����-���e�}�}dC��J�iΐIn�P[�>3\�B��`>��)쁬���m=�꽆v�¤�����Lw6�I�22����~�
k�	wy��@���W���T[�٨%�4�~�Z�.L�U=�7n�5^6ī�)�;��<�ߡ_�YN<�3@*@���T.���@�� �sD��P�{5L�\��1X� ��j��Cޯ�`_�ַG�~�I�#|����W��.2�P�r�)�as0�K���P`x6�׏�'ÁPNV�ܣ���`��閹�p�M�q�����D�w�a֣;���ȹ[�o���V��\Yz���׼�*���������d�Y0�������ʅ˱p�J�0jLMX ������xC�\��s���팵�+qqoF^s�Ɗ�J�rxF�H����9�2Q2���O$&i�3n�_�t|^��x���ګ�}�c#$�����8l�\E��\#����N��:FHs�+V"�LEְ�Lv4-9I[F���aȃ���S~eTƵ�Lm���
笾/*J�7��b91���c��N�m��.�(�5fY�����_��~
��	Aig����5 \�l惟(�"���$=��\lz�V޽���6J�������u�5�D7�}ҷ��R���7\!�J}��.��?��^r��h>��{L�����Û��E"�qt*_�W�;\�9����@��ǧ,J��#]�%Lt��JV~uq��sG`�iZ�8��"}Q& ��N�Y�z�/��(������<Ę� �;]�=km9a�mͭ(,P�}������+w,ff��y%8�a��Χ��h�����#s37(OYg~mH'���hg�x2��`N<0,˯��1��������^c�'��<*Л�a����j��"`����Kh��ߌ���l!����GU�	�}lիJhI�B�z�͡P�Pm�mŜ��k�	Z^���6��K�[��v�	�C��O6ZxGh&�
��yE������ ��4�u�;>;w�+q� "�GT��&�_.N�o?�r�}rw��|�[Ωs�aO]#��RJO�"j����x\����4�U�R�^�E���,�|3Y�O]�~xF�ɁG�d; ��{hs��kI�)&�ǀ�7��|�����'~�b�o;q��蒖�FX!0|ɨXOB�v�nƒ�ޞV�_e�O���j{� u��.7��{���x�Y1�:>G��Y��W�8�L� 0�fbK{�}��`��K[�g�:T��/3?�)��(�N�2F��}G�E�kW`�(���!�����DC%ۧ�/)L3��@X���Q�R�GV��������s��0�ʎ���2)�J�
'/Y&�orzG#z�P�Bq��l/����λ�9^�3l*�=ft{�>.��=0��;��M7�e��cnG�qa�)˵[\��l:�g0�]'�������>�o�i���<����-8 [[�U��J��
�u��i�+&q�vĿ��Z�6Fˡ��n�irWG8���ҕ�a�rhG��8��� ha$#K�Sۦ�}�Õ1��`����߸���F���jJ�K���o�K�ő�Vݣ�Vf�&�0;$��`��\#ʰ���a�P�Y@�u�\����E�Vx�/��f뼩�G����!�T`�@��0�&����gl��˟/��G�A"/��,�����K�a2�I����'}�6Ɠ��(�2\g��J$hl�+O�d���+D�c�Q���ҷ4�?0piTa��2�ob�.���˴���y����xC�ju�&����*�Y{:vF�?k�F68@\\�;F�foJ�\�i�AѢw�,�,=V.P����׋cs�gr�_������k�D~��H�d4]t��z���0����3��E�O����KQTlb'w��#!j��k�F��>zp-��WD�rfc9N���k�
�
����`)��Df����������)��]H�8C���n��i�Q��I� Rd:�_�0��*E"z4z[�(��/p��i�[��1��8g��X)h��>�ɐ����ʒM��@F�/���y��l���?����_(H!�x��UP&s}���9��~?��ey�L����I���ڪi~X�QHF������m�i�K�����Q�	� ���ه�6�um�#�s��_,�h�p�A�7z�C�+���o�����-P��2���k��%1�Dc���~���ժ?C��L��%9wxIcV�T.��̢�k��5C&�@������C����i�����q�2��B���Y^��k.�?	�(�������z�(�	VLH�.#��� /kw�D�����o���V+|������g�8-��5����\fq��')>��L���,7q�32lU����LW�w�Ĥ.|���@TIW<t]��F�!�[Ne��I�'�����E�I��Ɠ���D�1}Sw����C�����U�����0x/ �F+��XG�����v����B!9H�u����L���MKF��fR�Χ���z��l,��+� o�b*�@{��-�(�:�H�f������Lu�3->_�Kا7G�h�~4�
�%0<U�3(J,&b�O�2��|�z��n�3*A���ظG$�>=\�=�OqB饞d�ሙ<g
C�&��T�Q��fG���Qr�����ǐ�̍c���x��T�v��s.�� ���=�n]0A=�aMwXǰK�+�W\?m������a+d�J�sBb�K���$�?�����ہ~B�=e4f��g�#IH�~'iY?G�*����/��6��l��ݖ��}r��☚ۤ�u����7��,������t?���܏I�O�x��Fē}��t�ܝG�����E�T�@i�rQ5%b�5(�M�=��'���xG=a<�xϿ¾�������ݿ�MCs��r��(C� ��WFl�������q<q1�A��ӚY^gZw���U�����@�na�*�0���I�����dΉA#�
=3^��7fK��D���c�g�IJ{ا�R�	��6��[9������->ZF='VfRi�s����L�{_�c}�:D�8�K�0���ei�h*���+{�9��G�en#,���Eq@�/��Z=j�Ŕ��V���3&��}��0`�\f�\T`)����2����i�[3~.��[9�M�H�<k� �5���/�kc,�zw�����������[7������+��]��0<�	gTmw�YRCeY��T�R��PS�o|��#w��'��n(r�|�m�F�gku������v Wx����0S��Vb��vo��
�ʪ�b?�f�9��Ą���A$��!�}8`x� \j/�Cg�{dty\N$̘h�ɳI����n>D%+�	�+t<�%p&�qs����.���X���-��ҸO�uP����W�n�$�e��U����s�ޗ8�f�����8lο1�J�ym=�(���E
&i����D^��0W!ZYy(~�&,�Ʋ&=���:���k2���� ^uhW�Ӡ�ٴ�:&�D.�#��PV�Z��{��4��gq��#Od��'v�>�Q'o���/�׶'�����xKqT�(R��}�n[����Z;d��bb�w+dk�g�G���P������/����p�J���G?�R���Q>�-q,��9����/���u���%̝/l 	�6e�X��c|��o�,�6j\�1�1�b� �yc(�
�B�zY]�\:Sx���ɥ�RX����Vz�Ƕ�J0�����NJ�"S�d�&��T����m�s�b�&.Z�0b5�X�7���~�wh�D�>��!x���^�G��3��,y��),F��h��	�-\���$čj�૵���9Y�X*ظa�7gO�NwŚ<�y�z��J���Ӵ1��:��F�����N@�u@�]9ᣪ�Pn7��7ط0�C��:�On|O	�e!Oh�5o|8-�6N�aM�yO̪ϰf����و)n���~��=Γ��l�S�t�xl�i�6[_q��*�57��$^�޷����l"�<r���!��9�Ich�F㷛
%�}��uD�F4iC!z;�ᩔ��Zm=��
h�}��$��-��]R��Z�V4Jn�i�D�[�Mb�ɸkgo���H0��}�\�(A��_����*�΅y&|ICb�dC��e�ܖT�M�7"SF+�T�]�D)O��b�X