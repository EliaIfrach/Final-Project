��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@Jo	"3��a�N��H�m�����̭ύ�%?�EuDY�`�5��md}M�'�\K܍l�5ʔ8���7�G��@���]��*�'���A�]��I���%�[�n�'��%a��m�����#s�
�#�?��C�zC�>��I���'㰷�I�L����&z$�6;��f:�|'�>����n���Z�{2!WD�,pF�>P+�ߎ��J/�x��
4,*0�&j����a�m=�2i�F=�3�S����|鵢��Z�E�1.Q����=�G9	�"��x~/��y	߮�X\�f5�2�܋<=�S���v1J���,mB���ma'���)�8���ÌrG}M�����adA���B��+�q�=uG��l��~��l�9' (��`i�'��ꞣ&�I��sֈ5�q�ctw.�k�7D�끸��(s�$���8�Xb�aX�M��oS�X�[��\���7�f��맹���SE"tTLK�6f���e�D]��(Y�'=\�;9��֤I�M>ϯ�׆3F��&�^�~h�B(;�ld��'˭����1T���IB��;�܏���4��i5���e �Gܔ>��见1�lߌ� p#�q��0�F�
T2��e�g^4�3�1V���ho_�aaȿ�^Q��|��\���F����F&�r��7K���s!����<R��Tg�;b��J3�Z�nW洞��x����Z�	�ܯXae[���tiä�g��r��$���ၵ"lA7��s�ٓ��Sy��(n��ډ��M����J�w�>�y�B2�{=@�&�����L����y ��Wb*E�p^C�����4�ȿ%!3o&H�i��A��
��x~�3+��s���)�Ba�$9�*p�W��Cr�Ec���ں�L_��qQ���N���?��\��L���b�7�&7Cჰ�|%@��t���Tp�P�2�N	'䜣����GG��� ���l�)E�I{?�@��Bm�DMx�{��J)����I�?2ʁ��QP��n�ȯ K����7M)�8`�&!��VP�|�mr�i��RNO �â��d�J��Z�c������3���f�p��� ��q(���J�h/�,���\uK���x{��'�
#�
!~t9�-.�0��GV6z���SV���N y����� ����������FR�?�����|���CU�.��v���g ��k�����ܱ��:6,=i
�8������+��y6�rw�~�{,�~d��i�9�ް�«��ʈ@H/�����ɤZm����?2���A<Xݰ ���ϣI�k�8����8>
�*���2E�gEH��+
-m��X#��^��
�\��A���E�����ݴݠ�,��^V��m�~�\H��M�_؛f��z��o��L��#|.͠5�|@��-|��o;c��A�OF�5P�2g�}��8�xj3����Q#4.���Qy4���˃��^���T��ς���[�qh~����]�;�� O�z�D���k�B�M������Z��pP�PX��J5*��Qv����9�U�M�{P#���yx6�{z�8� !���Q�U�=�s��t��!X*
$2~��ӑϬ��N�7F�]�oZ.Oܞ����p_��~y��*~Y���F�kat���B����2���x�<�)3 ���~Kg�.�Ye������E>�V������" �YW�!+��m�r+#���ƃ�AB�_��	D��<av"O�yL�Ѕ
�Ӵ;���4m�2��q~��6G�P# a����&i_]�sZ���]y����c�xF&�J@lhpf�͸���� �����Zx����Tq�E�6����%OX�w���z-�>b.�	�z��x�gHR<��~n��|�^K��{�ׯ3vsb5D����ނ��E�m�˯"M��9�l�x䬨�?n�'�Z� ���jT�0��JU5�?�ܯ%>mH�>����zl_Z���i�~B�����v��[S�d&�&$bK����ɥH,S��.��ʚ��)A����V�f$�4e�U5]d�7��UK9��eO�r��_Z��Vʪ��,�|�<w8�x%%��0��P�֝5e�D�]�PX��2f�Jٚȱ/KW=�rꎺ���IR�'<PL�pZ�B@%ג�G���i�C����,����XX������z|�4v��G�>�+dXy���\