-- PLL.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL is
	port (
		clk_clk                      : in  std_logic := '0'; --                      clk.clk
		fifo_clk_pll_0_outclk1_clk   : out std_logic;        --   fifo_clk_pll_0_outclk1.clk
		reset_reset_n                : in  std_logic := '0'; --                    reset.reset_n
		system_clk_pll_0_outclk0_clk : out std_logic         -- system_clk_pll_0_outclk0.clk
	);
end entity PLL;

architecture rtl of PLL is
	component PLL_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component PLL_pll_0;

	signal reset_reset_n_ports_inv : std_logic; -- reset_reset_n:inv -> pll_0:rst

begin

	pll_0 : component PLL_pll_0
		port map (
			refclk   => clk_clk,                      --  refclk.clk
			rst      => reset_reset_n_ports_inv,      --   reset.reset
			outclk_0 => system_clk_pll_0_outclk0_clk, -- outclk0.clk
			outclk_1 => fifo_clk_pll_0_outclk1_clk,   -- outclk1.clk
			locked   => open                          -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of PLL
