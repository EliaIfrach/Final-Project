��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
|*�\�MjC0zP�����^{���N�<N}@lS�h����C-6�[߾&�9�*w�(�寚n1W���a,����0��k�㎝5��X�ҫ"�лW�㊯�{�Ym��^�u'd���u)�DC饅�@��a�\���\^?W�J�HT�?,o�!u�q�͙�=���Z�cZ�4g�r�K.-�jJ�Z��a4F�?/Z.�ؽl$;_����>)_���1�,�6u9s�K�;�������T���Ç�5���;jC�Q�mzv���g����Ȫ&G�t��D3��(h�&:aL�,j�o�h$]^	ky�c��Hm!�ľn���ʶ���$+��΄�Hy;���\��E*�. G5���ŔYd� �<@����9��.��gDd=�����J��nY
l���<8{���QC3�����{�No8|c�(�����4n�����N��[P3��4�ﱇ�1����~��-�&K�4�ӂ4�f��$��Ng��¦͍+Ύ%����q�O'�0�;-�K\0LQMMkX�V���|�;C�(�*��/��1&e��(r����������+K��	���a��;JS��/ݯK(�
;�Gl&=q�f	=��ތ�M��K�9�j$����\1�<
#��
��k�j�}l1�<;�臄���*> �����盧��>o�|V6��Io�K��+�=�����4���Oo!Tv�b�����(����eca!
��.3�������Id�rA��;�0=i�w�� G:��Ѳ-,߈O�G�#���<u�[�,����ٯ`d/�	/���$͘�w��EQǦ�~�mc�D*L=\�?)���	���k:<�����i�wS=�����Bp�A�����rȟ��ӎ�0
��f���@����W5��D����v�lI�������\����X4�	V��)�/u���%m�Ʒ�ŀ�7����g��ͯ%�1:���7�q[�ZX������e1��6��	��n	�U*�-Xs1mw� �k��)�չӷ�e;{�Ґ����+I�O�4����.�4�H�2���~���!|��z������C_TM��lb4�Ǎ#��#i�6�8@ߕF��O�p�3$�H��l(�э0��Sx���Gk؄>fC�] �^����*���!��1c�M�-����������t�&g���mggS�`�$8 ��9$I:Osg_��L����
�k����~��'_GQ
 T��Tɨ:�)*epa,`�r�ƁOD���O�mETxII�2�o+x�N&��X���L	�i��v�������gK2\֪NQf���щ�n��={<�����-�]U��U2� W<�3���$+jA�;��,�#8b"мM��5�3/gl����{T ���bYO-�Exh&(�o�����bTe��EfO1�GU���mV{�GeB׳p��<AW��AxWHH�	6,�������A�`he�9�qn!�,�(�i��N���6s.�6��>ڠ�����_T�ݦ��@����z�ܴ����m����S"�Ț�		Cx@�1q
��@�������;l'�HY���l���}ި-+ۼʏ�ߞ)��u?�-ʹVy���Vu���n����~�k���\�O�#c�1�)?�Q�G�D1H��V�EV+��gݎC�0��|�RV�)!��.�X��Xp[|~���J�#L����{�8���j�%}��� a���9=��hi}�%BL�8v�ʏ?+�1A�A�a�=��	e��
:���7Y)�]�R&vě(���4s�FQ��j�ꯅ��B �Y�'�o>��:Q��k�r	�P�(P�(>j����9u��p�Jׂ0Ð~���nmZ�p:�x��r�O�!6~�4�n06��ז���v?N�Qԟ]B�p�m�4W�R&,1>'�ɑY��5��5)QaY�9ZFT	~��VLq7�=���X#Y^�'Lb �wA��+Fgy�<Q��C�;��L����6�
�J�S�b Q�������b�\�-�Lܙ�W�y 5l�%�y(��k���&��zǇ}����>�-�`p�Ns��ĺӮO��0q	�%�h1���TlR��_C��kc����-�tHd%s�/���Zq�咠ع��{�����W
�I�ViTƔ!�0A� ��&�Ւ�������v�mJ3�$LѲ�7�y���i�Kϕͤ��a;�h(s(f����^�dFE�x��w+���W�&��peU���m%�]�f��\CĄ�Ex�b��ܣ�xr�TVN��%� �6/�P���8��栘��d�r^8�Gh�1��L%?�e����+�$e�}��
�*l<أ5g�\��j4�<��h����2>΄�ڜZ��v�<��c	�M��({'u��6�/A3A�5����OW��H���s�ә9�7�jM�a�}�O�����U9m(UV�V�ndc�,{$��ԃA?���q�r՛�Z�6�A���^���C �B6��ل�d���K�3���N�y �r��gZ�ʳY�p�%�ٳ���/7x�i@�"� ���Ý����s��"�;���.�ug����'H�=c=Y)�b̷�C�i@_vQ߽�d}/o[돿p}����i4��Lr_ף�y�K�,��L]ñ�ij颥��{cX��2L m���D��;�-��t�d�Oy$�����	^��E~�ao�Ro�+.�Yeq[yrlJ���1zM��f>��SbO��_oc��*�齯5]���Ő�Y�l㻏��3V�f_h�ۇ�lIl�������D�p?�Ӟ�A�a:Y'�ǂ)�ѻ�z�<(PNp�ᢼ �2�7�&K�&�f����60#EZ=!G4ن������[�D{��|\h�,92D��+�/h+`I�U��Z��Z���	�n���3�q0fd`�u�BǅY�:��M+�`r@���QG��H�:���%�c���9�^�mYb�?�a�}�C��~�x�f��B��7m
��Z��V\����[��P<G��0���ťr+�߲,D=�y��b
 �*�\J;\c�ʵ��v$Uؽv(�?R1�<��]�&�"�'��ɘ��3a�˹��C��J��E�ì�))����N?���A3���N��wb=p�)x@��ZV�|$��ӂ��\�
 h�k�r�Ԭ�$\����K� �L�Ò-v?$�bZ�7mI����W���#�єK�_����Ӹ\G�c[5nN��ݱ�(E/ay<��P�oRmJ���â� ����n�Ed�]1eҀ����+�a�����g�	Z}1�ޫ� ��7��{D����غ/>�\s_�����ju�$b����MQ��j�B�x������3\5���H	����ՠ�y����!l	�V~���ɏ���P)]#+)�E�u,&t���O�bt���]U'��FML�fGD�Z��,hN(_R��`��qQh3�b�����" ��̌Mn���Dgw�I[)�L��sm��E<Oe9��
�K�P�ea��Ym�5t��#���ƨ�IG�:t{E0e1���q�Q(y��8�dS��o��i���Fq�c�~���	���1�Ej����L.*�f+�D�>N���I_$�E0��k��2���Q�¯�AR��|���ݿ���u�!�zM�D��p�&W�aב>c���N �kPC;��=�")G��!=�Lo���o�²�x�;��c����s��,6�y�3Y�+�ʵ�̭A�#6�����p���G�m�e�&����&�$L���|�f�
Hd�\�ᜩn_����l�l�LAQ:�_�k���ݼgĶ�u@H�-���A����%���(�� H��Tl+fG����
ғ�ȏ�	����Aw�zz�G�$/�n�yE�hr���F�����Q��!���\�g���H��+��@Z�5�r"���Ri
.�%�A��ZG.|x�v�ݾ���NL5�8�)�ű�Ն�T��h��֓M��1~X��e��qx���J�n�!�� $[G��Ҷ��	x�t�����$X���P�N�q���ƙP�K���nΛ�1����$��WΎD�2mé�f]�T"�̶�P"�w�����z�M��D�4>�Z�"�p.�3|n�!��)F��e`q!c������&ׂ�š��:,����q���U ͽA�;��Ey����m�!Sy 𢡊�Nͭ���b{�b�SU.l��[��.�я2p�3-d=�d����ȃv^��C71;x�9F��2F���7b�BGz��\�u�>V�/=�����9�}�[��B�i ���)�B��!�Q�{�@0�"��J,SE�Ӫ�)�x�{]n3Z�B��nx��_6��9Hȗy��&��i6n���������up`p��H��ř	]ֵ<X�+d�M^4zel�������7����E�����f�Z�[����z��0���M1��ʹq��F~ ax>���ߕ�y�B|�=�&Z�0T�I�+��t �㳘���ƌBک��=��d1�u���u�Q�DE�=ks#��=����Z�o�
:H�cUsڤ�:���yK�:y�<qE�G�?���4`�)v�\Si�K�ny�X��o��@Ϸ�����@��B�<�x[r[�R�j����~*�hf��i����%uO��F�I��P�+��8w�Q��/��������fM�`�J����y	g�p�.7�:�!և����ǙiK�4 U��+��A�Kw�m���T�zy-jb �I3�H�	��'l?Ӡ���`kl��duN)�s("u�'�Xi�t��������@�{Af�隆k6�C�p��}�	u���/+��:%n.&xY�������G���aε�6-�b�D�_l�I��Jf� ��;=���7��bր�A�*��Z>/��l\�S=&�"��e�q���A
U�sX?.Dsj��j+�D�R�3�1�Q)��x"%ҩh�/ȲdHv�xy̠6]3\����LQ�N�;����7wO)*F�#����2z��]x�U�n�у�'Ʀ,,;�db�UV�·��\���CL6$�樞G�jϼ�\���3�F���@l����R/v�^s�1�Éf����n���VUFk��]n1Bm�g6�@P�I��@?w�A��!l�07���A㎘�]きr��8�VV�VVD��l�i�).`���dW�K F �x�Ⱦ;Чis�W��_b;
��Q�]�.C��gcZ��ڍܼ��	z �a6�����M���q~��GPZ��7o�!fQYn��)����
uΐ+��V����Xu�V7P�GAE�]���)T��|��sƈ>����9	��B-b���ϵ4�D�C�d9��>t���AG��$( �!���6kO�(��ɠ:��(y�K���4���Pη	9�x���<�W��)?���}s�]@�Jl6ⵑ&�.cW���39�>��j ����{�m���}*�&ܯ�u��y��M]�(��m��f"�J�)�$Y��)��1.
Yg��<��mf�Ө96hW^�Vɚ3��ZJz�������3ձNz�hoC�d~���Y�U{~s�8N2%=<w5�Zsy�qs��S�9G���.��p��ӌK��|I;q������a�W�t�p�X������ޢ�I#��)�\�23R�\�,g9���x�c�Mly&�>�<�G	�/��D��Ue����՟p�r��%��AȪ��W�v��+˧�!&��-��U�4;�j<��B����	|/?�}�30'��`I��{����z�BL&#�������~�QZ7�Tj���E&w��.W�l��η4�KP��b��$vV
C���/��A�)��[;!�Y��{l(P9[��W-�����#��4b�����;mMgf����t�1�k@ԇ�Nc=��r\��8-]	CN�B�Is甽,�̷R�&lQ��Tx�d�g_��"b*!�򲅥 Ҽ>�ۗc�W�;��~�h7��g�R�d[A>��Ѹ���}a�]��M-x:V���\��
F���K�)@z�X��E�QBtPuu'X耤�v5_��G]"����w.�@$6��
��z`���!	l�Y��iw=T��4���F�$6^9���,C��lȩƶ�	�ؑ��q.�$V���%�7�)E����1N`�?��@�}4Y+���UӶV�:�Ԅ`Z6�y(d��I'�H��a��]���EMR�P���j	������i����� 6)�;a)怇����$��� �A$��{��^4�1|r�.�iL��+C�<;�z�Q~�Fg*lP
����?�;~�d?��ذ��ۡ��8 �Kl@�g��e�O���P�2rwƾ���A$>��<�o��>��ѧ�qV��Y
������,b����=���ˤ =3^6���5�K�"�'=I$�:e4/u89�TZG	�Ő��G2m̷0���[����,� B�ם�r�1�|{�p�w�l[|�����Ee����H�?�4K�
�\�Oʞ6dY8�
c�4S&��'�.]D�T�:c�"���#�������G�W�g���ۣH�� ��͏�Mz�׸��c��Qi��{���VG��؈�v:/���Bjh�Hg����������o���� 6x��ۃ( �?�����>Ω�n�=�_%�Jr��~RF�.xz�N7ar������
n���xˮ �<����tf.�B�U����� �\�)��';|=]$Ũ�	���qȂ�(r6^E�h�JI ���-��(	FxHa�X�����& �w�"<@� p���&�P�uڞv�J�%���j*�#��Z�?�}��a�L 5��N�*dC�����ǫPw�3`U����+�z�j^o��"��8{I���'���p	�_�f���W�B;��Ʃ��>��F�Іet$.����F�F�ye��`j�Q�s>�d|aA䊣���7��n}M����>"�f����	cx�AvP�5���y{4�D�+]�xd᭲�&���{���(鰇�z���QDݛ~�7����ϒ����� $K�5�NH�+����e�票r��Sv&y��Egvm6?���[	h,�%�[�}!�e���=pyڒ#� y�łw���syv<knR���r���lq��E���@�4�������� ��������j@Z]WE�?�{�[������̼����0;����;�Ÿ�@���u;�M�"�fw(97~RO�|irY�y(�|zh�(n k��+.I)Q� t�{���g��Fs� K�2.���Wi--�F�ڣ�'��$Wr�;�"O�hǎ}�Fo�Վ�f�:C&`��}��$��� ��:���UA�:��N���^k�]]q�E���/d��||����c��J-��$�>��c�{X��dd7�w�+gQe�����<������l�Mn(��"��)%B�w;���{��d�X������4�:G���O��I��S`�z������w�(ؐV����S��d�L�x�wdjXf�=��i~�o�+�%��q2yM�vZ��X�O-�e���7�s��p{*�x�����b���Y�|H"˳4Q�X&�J$��	�zz� �}����F;��!XS��x�`޳����47=��������rY�F�;��QQ��cѡzC��ZQ��?7�)B�
��G�N��O���T(~Eg0�-�Z�:�sV�	�GtC������ك��k��Zn����&|?jA ��%xV !ގZ�D�n����G�s�6�*m�B����-pf�+F�]h�Q�
's�hd����72��^���ME��:,ɌW�P��jQD4�7���ˌ|��մ]��ڋ�7������<]m�']��^�^�#�z
/��@�l_��;���^�jK�Ȝ�_���D��"��Z'��bo�-�O5\� r8	�؁��8�6�~�vhQ�Aǿ�$,� �c<��6.o�e����p���s�#���fk�]�nroje�����������,I ~a�����0�dQ�d.
?Od�O^�89���Jg٢�4���Ef������}��k��rX�R�}��l�k��!��l;�:/Aa�\/}�a����C������!i�r-�n�>K�8�X94�T}�L�[�<�/���.=�E0U�vmŮ�����>xu�y��SU���ǌ蔙y�����=��B+f��#��/�~��۶!iZ0��D���'��j �Q7nN�M�|EG��Ka�Kƍ�Y�6@p�>|뗤1�����k�7̎����I@��-k��C�?�@Q%m�t���gj�u��G��s`�K�,�ʛ��mU�g�c��� �|�֮�>�\�:ڦ�D�2����}����B�tR�ؖw���9�91��P�Z.� 3yJ/+��~,��N���ٵ�6�|��(���H|���}�#��.�0�I}0�h�N�;���-�q`z�|`��^γ��r��ff�QĝF^���)��+Zt_sQPX���HKd����.�������!_�^N��'v�K�M��6N]����i�G�7�]a�`���BwT��F'�5�EjoH}zJ��٭��)�u��˄�L@����W��p��~�s�.�t�5��#"Z=\��ө�VFӏ�,sw-?���y��6Cx�t��#�n���A��;~LY�>�f���k9Ks�haĿ;��ߘ����`�������� ��?�\@��p/��.�%WXJ|�<���؈1�F���B��:�Ib��Q�S1�s%��ܳ�6�`��lN^'�e�~�h8�`u��~pdYߢ���w���]Wl*-��Q�()���:$g�}��pq�墱��e���K@�n�A���fj�^˂d-��<�l�|�NC�ܜq�)�$.�g0��N'%3���wؽ�(�� �U��餷�,S��B�J��,� k=Ge!��:�E��7�u��4�,��ŽU��opD��J+'�	3^!�M2~c>�q�xO7�ʚݑN��A�2H��`4��X��o��,��"�A�����{�w+@Z�G�θ�7%�����4�����j&��=�#+�WB���T(*,(�����R
�s�BQ�Z&B��$��_�����{`2���LLnr�a�x+PL���"������x� �6��X���_�@�\�5������G��F9��^��A����VUV�,�y��� b�ch�q�O�2!�����|�MC�d�sx�$��*g��mˠ���n~��x��1ˤ̞�낮Bf�ҽx�M�+�.p����(��,�r�������X�}�6E����1������q1����cı��f�<a�o�����m۴��� �ǰ_D�ބ�)]��a��s'58ԭq� ��*0y/�%�-Jj�ÒP�r#^ �	c��2��
�[!�q�M_��FĻ���?�W��s%O�����W�����_���[8 I�A1p��M�?l��)%~\ݘ*؍:9=��������v�I��﬎������9��r^
rTE�.�
�օ���ٺ0��
0�F�F����b�d���ęQ���0����h�g�hdF6zП�l����2��
1�q��^��q*��\�u�G Vc������Ds3�_L`��.��0{Fj�Ʈ���w��ʂk��{2/��7`�����!&�_r %Z�㐫и�Yj�>ͥ;��^�������G��ޞ�����N ���+�j��H��������ϖu�!F;�b�(�W^LP��Q�A�:RFϨ�^�ߨDmE�oe7_%%�0*",Լ�d�L�+���m�{�[E�|��C9�8iÚ􁎳��^f���?~��zm�)t��e4�S���[r��������;�nv2��w�RP�5������/ˍM��K&�n�P.���U{c.@�t-@������۔�8��I�}ްMjr҂!�����V�����2>�j�>#r]�c��ԣ��o�V�-%.�[1c&/y��U��%,��I.�A<$�����)�}R#����X�S����h�ֆߖ��[ �.`~�vv�l�l}10{�Y�y��4���C�sW1hE�����]�I?Q󎨛uݥRvF��KSI�9�����)L����@�q�,���%����nW=A��D/�?�������yix���9��@��̴�����Ur�.I�ʿx.D�"��L��[�-�m�1���܄�����%�s��z�()�=�ڈ�(m��~�����Z8ώჄ���tbt�3����t���/e8�Ϛ({B�O�9ѯ,H��i��a���:��'9��Ͷ��_���m��~�`�Y�����l�&��7s���œm�Y+�V�E�Q{}�h�QU���p�႖�I%#1 t]��=/e��n9���5VD�w�RY}BMw}�hbB�"�Z�ϥ��N��t� ���U�g"�e��+/!��uJW�'��ҕ̘�^���g�c�a�H� �	�qSfT��H����]�e��=�y�<"^�mNc;Hѻ�8��K��;{�빑���і�\�H�����i)PO�����$�gA��
��m��/�c��)LT�U�GSF\�ddFi'�%�OL����1�����2���� ����a����uy��~菻�����[�49�tf�PM��PO�|��g}B�1y�5��K��5v��:��"����;���p�����0u��jQޤ�K���4=IG �%�����EsKm�k��Z����I����;����9+���33*9�t�E�=��]>��ϸ����ߑ��}���%F3�[.[�;P�ƽZ+�u��Z���a�6E����A7��U��'���s7�g��7I� �ygs�X�hl�	���0� ��d(C�	�P٦~��Xzc���r�(�k޿�A�,�H�R ��h���
g�Ԅ�+�Qw(ꠃ���N "�>e�ŷQ.�4�d�2~v��h��$g��n��W��̏��od�u��lE�m3��!,Gf$ %I~j�t�z.��~Q�+�)qt�-�x*Q�Y|�X�����$���Q�oܣC73��Xɑ:�=_E����b������� `x���[���C��:�3o��V?�~If���|�����*6@k��;�����F-��b&�
�c�a�~���-����&�o�lF
����-�6w�*�Z��\� ���������B/��<�����X*��ŕ+AÑˏ���4��G�G`�5�@��Ͻ�8_,���/�L���O+V^o�P|b�'�0k0�M<2����Vf+@<�p�R����R���|?��Ooo�r�R�9�X5EQmZ�j$��r�����1�U��N�6q��O�Y X���� )�ٜ��n�1���#Q�|x�͒_{G̡��OϽd���3�Op�����!��$��5�e�bcS�wV(�*Z�Z9͇��Ot����B��hϥ�/�L�������t�ܲE�890��.��*�D�wM�wu�գ�V�7Ȁ��V@�9"�XLZ�J�����:����3c5#0Rb%��*����(����B@Q�9�	���dY�1� �?5[�J�Qp^}D����&�	�ɛ����]>��WY�w~���R�k����yi���>z=?��Fbl}�&,��a�x(�fE���� ���_d�8ܭ��ncS�mǋ�ܬ=�UP���[K���+)vC3fCԃ��n�\TX��$hNN��N��������|qu��k]D\A�p�]{"�s����j�l��J�~,`��AJn�7e�Ѻc�o�O���ի����ev���6va�ֲ�!��uA�,�������x��te�g��̺��u���`t[6�&�?ڬfv�0�ם�� �r�y}l����pؐˈ�|�WS��q
�5"����EK�0�}o|�F��p���3:�S���1հp������\v�qe:u�:t�4\u�^�Ք�1lܬoIQ��ML� ��´�R�"hu��xp��s�|��j��dX�+RT%y1�ǡ|�����vױ�W&i��V�PSR�x7�q�`&�L�#�o�AG�Tp���d8��izl��o�9�!�LN?�@@�:�w����%hY5&}��kA�K!�58�6�9��
�缝������Qp�9vKh��nL�����&���4+�@q��r�yX�n�_PHɈ�QI�2�O��$�ž��4]Y!:B��j�,U΂�EA���[v%ءB���9���l^{��ceU���L��i�c�s.�е�KX�GF<�
�t��R�꿎 Đ�=�oU��
|{����%��W�ۆ�*��+Tl��X�R��k/�>�ǵqUEdźNY�x ==ܲs�qB7�1�80��%��IwI��Z`# ���m��M�(��P�Ao��� �Nw�/71���C`ki����5�"d��Dl�D�Z>K�Nl�%-,8]�-��E��S�	�����Yh�yzoM �~��m:���83�6��*�i���!��m�B\� ��Q) �
=��UQa�o�<��oG���	쵰3��\��(�_&j ��p�Ri)@���1@"q�:1o�5�:|�ۯa�]49?0}����ʂPrP�L�f���e3�F�/"2�(F�
�s��gp���e�JEs���@�A�	��hϛZ���'=�y��&P\�m*4� �,v���{����hU�\V
�Eƚ����]�v�5�kv%#x
�I�5�!O���QG���th*��ҷZ2�{7>s�LD���G�$��/"�{*����nS���ʜ�Kj/�|��_ �JmŜ��hp�L{>������p�%Sc]�P�N�b)2{�|�%��+E����w�޾��I�H�"h/��$�H����*����kQ
�$U(��J ��E�`	�II�!o�?�_�=.o�@]QH$��A醁���&��{A�O����_@Ou����Gw�D�mL� �>�I-��g,����OdG����������'4X����SؚH5&OO����p5�i��:��?�TD��.�t�`��.z��픯����"q�q���95���zNl��(K�9Px��aV-���!��g<,.g
�y�8=�9!f	$�nZb�=�R�@�7�5G�-GVrB�*x�/
��,(��I��΂kO�D�CT�رI�N�85Z�H�x�� v[���%�(�%����:�kA�l�<G|E�;a0΄�.���BT��>��WT��i��S�YM������ E��9�g�C�� |J5y�$B��{�WX�?Kz��܁��G�Dc�>��HRL=�����e� �vv(d�6��67���}��e?��&�Dy��V�W��f��^=.�`��h�_���R�x���։hft;��*��E2+c ��%����F*54�wYJ�<�һYd��ۈv��B�����/%�-�P=cH�����23��3v��Kei5��2S9�Z���f�m<sԄ���;It�S'��	�=sޫ�����iGs�Ϡ���� c������8��H�K��k�E���:�Gm��E��"�z&�sp�Vp��v.�2��
�Bi�7}��wK���"���Lf����p�Sz~y���>y�<UW�r��}_��m�{�-���F�s}�/�e!���̩/�)/�iS�HO$_�ν�
�!�HӤ=9fX�?�E�\����@1 \�O�=�M/��=Ѐ�ƼƩ��M7e�	o3���e�r0�yo���H����H+�5q�;R+M�]i��<�,��j�`�ҥ�b�U�h�S��f��-�i�`F?�H�^�`���_5���^���*�>h�B����	�LgW�<�	lP`����J��5*E�apC�ZX0l��]�m��ͷo�N�1�"�M�{fߎ����H��|�Z�1�;Us���A�tH��y4������gr�N���y+��WW%��H5�t�|0H"�� �2@�����s�D���O��I�<0��q�_�kֆ���)WvD�.�Vz�E$l�d!$���	�1n�-!1	�b�k�I�gY�YWr%��?
���(�H-��rp��Km%ǐ��|rt�l���ﳱRƥc��X	P	���#�˲'t�34�����U̝�e	��G��$���(;��S�8Fpܛ�|�QI��ib/�xG�i�DQ��9D�B����'N@K�sp��U!%��l��mi�}�I	�*ܝ ���l/]<K��Q���rvu�o��ZE��s��E��5T.˺�JQ�LAd���:*���4��Pܶ�v�b��+�wU6���6lNr�*xy�T&-g��Z��ܖ�zsnoG��~�)�2��*�j�_ɭ�M��dJ��W������V1�':�:�a���^��_��`�>���ǝ�7kC��A�|3���]�{=|��t�;��xQH:�͗���!�/�aAb��4����)�~x0R}7�ϸy�uZ��6��u�T̆A* ����.�A����9��*oZ��R�B.���I�Ƽf�M��n�͌�r�jd�6��C��c�/$΍U���^��Y�U��Y-��?���ܮ�3��-+��T�5�>]!����&L_�y6ᇳ'����A��*<�]^k�����§��3�X؜���l�]h���db���ۼ�!���^���^�Y�e��M:?����!8��3-�Mi��-s��N�!���*��)$g/!a�/�����'��*k�ڂse��⯗O=�Z����>R��xb=���Na3 �.��玞���� ��`�:5�@#aIs�k�g��-$�-��\	bs���)9�Nٰ���w!(aHP3:�;�"c�/ ������#�H`Q$U;O�Cp��zHc��6�
K��I�oF��Ωvu/7w�i'T�V�P�#o<�e�b���b�O�U �<�J[��C�Tt�5fOYr��|g����Z�	�SP�����l�+�"�<��d��ݩ�S�.٘ѽw|�� ��^�k)pI��8J2���?y:���Ҁ(-���'i,:yf+W���lnz�B�4��ż�Dz�k�L��\��]�ky3�4]C������V�DO��a����$����yM4`\5c���*��FD���xz�*^t�|����?�"�]� 8^�M-R�Q$c/<�� ���x�y��ż�A�� gMt�orN�{e��GYҺJu*y/���iK�v� �0V���[Yg0h�2�-y��AvgC��z��4 *s8�m�1s�
"���27��w�Ss��A�l�Thk��0����Z�v	u����c	N;�W�F2�T�K�4֢>�s}y5u�	�`��n���-ip%1+���������ٝ��S�d�C�Zت�0����F��8�l�3w?���c}È��8�����ط�/�*�BD�B�/�Q�8cf����͝m�-�7��YQ�s�����1�����d#3�m�d�SJ'��~7,����Cn���/�������	��6�?aS��W�*�[��{�wu�gp�ۑ�\@��`��\���֮&�\B+�vBJ\(g�C!�j��N�.�Р�L)դt�XM8v�]K��TC�̐�� w�#+�*���~Ňam#0�E�Y9rC�H���|�8� �5��&wVs�\�$�n5w�ea8����8x���fؓ��b0���!G{v����)k�d�)���]1=�zj7k��Jt���ך;�?fRO��C��BvFo��'���� +Tk��5< �D4���iSb��e�z%D�_��W�Y�l:O��B��:
�B�&A�1kGB^́���<���-���J,����8�P{�	��UXg����Փ�Aӝe����*���)��3U����	�m��2��N�SC��R�E����Y�&�=�s����=�~
���U��M�H���ɱF3�M�����j�k`���m!D2;�ɋ5���������nW� bJٖ�pM��`e������e��UW|��oU�XkK��k��Ex1�ɜ��̩Op�F� p������V��v��)R<|7� B��o�U�X��
�A|hJ�Ѭ?k��g<���:���e�������67,mp�;�#���T��y�ב�#�PH�ʆ�ï�i6{� P�K�Ӥ���V���c����[�2� ޶�Sq\�l4�ؑ��$}���u�I9����`d����8�x��r����q�������&
l���ɔV�V ��}��C`�i����%y/�AD��YX�Y�R����ZH��C��e�d�1�E	������Q���ݦ��5Q�Y���q��М��[D�x>�s��M&�=9A��D��a�W�&'�b��|6>;��B��n��a���]'��kC�P��(�mb��Ӻ1K4e6�\��H�j�9
e��2����>��b�]�2��	9�<�b�r��ňFL�39֝_�,o'���.?^�m#��UvQ!��x���Vлu;�\{�_/�����7i���н���l�_�0mh�*��z�T�Hkf�&���s��|��d�#���Σ���yN7��g�XNB�# =��VM��.C+ 4�J>^����Ǆ[-�j5"5��7��繄-�)N�����
�
/9�4A�Y�,���I�(]n��� B;��C~�1�?��?vxG���
'�9@����<�)ce� ����>I�G ��Q�>o�����U�h���V2��72�Ux�19�/�!<����z��?�r���9�ߐ��&6�t)�TǢ�7�� M]�ҫ�j�i����U�k��|=�:lu��� 3gl��@�W��gP �F!uN�4�_�\o�h��c��jH�kg�?�?�1'PYO��(b�jsu����TE�ԅ�Ⱥ�b��¼� ����W�7˜��Y��{^�s��믠u�~Aqn�}m{�.��X�2^�diL�w��_>,+	�#��a�^��v�!T�x,�B�Q�����Y6دgS�`c�m����U|\�oD3��~�#�!fa���3Ϲ��
���X}:�b
���]���m��X�ZMJ��>Y5�65�L��W�cz(�H�0�~��L�O��6��}�QfØ^-��~�j��O0_;�������54ֽ�vqk��,Hb���P��M���L�V,��!�t1�5�`�kحI��� �{Z��D� ���|�ί0��鳴�����dr��]֥\����������~3���#�G�Q��:*SZ��aR��lo+d����T����멤�DJ``s2c�, �lMig��ς*��2[�q��v�����:IB�gC�7�f:����O����\R/�
�5�nC�]�spP�������T��8�S���c��KV�*��)ɪ��=�e)u�2���v��r�C |�^���$��WhMѷD�]�0*֎��)��.����etq�1A��o���̅*��OX�8̗��V!�t�6Ox�f�y�;��ua4�e,�
/�L˜s(N3S�M�bjJ*�k1O�V�f2Y��Ӽ��-u@�i�.�Lr����!4�g������"���Z;�c���SBB��ˈ5����iW!&��6����4?:;���'����f����Ua��ޛ���G�B������c�Ge��	�j�ͨF�����N*��td<e����x�[T���\��;-����`l�ܹ5y��#��i'b���(�^Z�{��7��/�0�Ā� A5���3�:",�M��3N�}n=��߉ms�C�r|dX�U�~�~��{:8�r�P���.����@袰l��R_)`�O�	��ɮ��������ugeGp&�XH��H<�k:1� D�r^�z�y6�&T�P�ۣ�9x�v&wN���,*㎥�H�ݯ��д�e��T+Je[VZ�z�"]���m�yÇ�?�٬z��͐��=����ѩ��#�S��ٮT�-������-��?�Q^��Yy��
�2[>�8�����!c|�E����n��bS��4:�ʈO����;���k
bL\ Qc����G���%���'G�Ώ�����<֟	�y�z��4�}���f�l���Tu��Mͧ7YJ��z����'��h��A`rh��%-ۜ�=埐cG��P���T�7.=�ʉ�TdЀ�3$��3���C��9|j}�&��R�!R��Q�}�
z��a6�E��J{���sR��!���*;Ɣ�c9�Nb
-���/eMI(�}���^��|Kj�<�G���<�A�Wǰ��}�B(�?�J.�k��Pf3IEO�:,繁G�Wu���d!�@07���^��ु��OAU.@� ���XWBҸ�����	ݝ�!�	ɷ3ԙ�d��OE�/�k�;y<ǈ�h�:�R[zUR3X ��m��a/tyb�W;�!���'v�#s���|�M��}�j����,�AaO%e�R��ܘ!���NoA����.����aT=
T��Xg�`�	R%�)>�$&�yr�roJ��,G���N;KRy�N�N��Hj�'Y�q������vN՘Lǯ �Z�Q�w�T��z�9:	j�/z������0.rq��,��5*����L�'���Q��7���8�h�:��	|�0���bڄ# LY�$bbgc��n~qy�jG�[O�����T5�,qO�j�8�E�|�w�`�3�`�}�7D^6��0R��ið��ފ�šZh�R��<�>��{��q��&�f�4o�it!�6�7�ג`��� h��D���UuA^��ep"%w�Kb��cڄ�/!�F�!~��ьwWpX��ڪz�3=i�M��>�1�{3|(X��0y4�F� �g�!~��x�ܶ�Sim�Y��_�̗�o.A���Y<�ě��A�5�e/�@m����O��g����t�c)�7�"ZO̳��<#�H�E�b�kM�gE�B�<S}�m����n�`AHUD�s	Dl/��c��F�S��+-�c�H��N�����=% �H=������h��+DB:�A�`���W81�	?��Ps���o�3�p^$;��B~V�.��̡�W�1�d7H�i��+����������m!U�g�� ü���3O�o���&���N
E��#^�>����3�bQ���� �:��M���8[�-吼�#A>��G�՘O�^[��>;�9Y��!x�Y0�ǔ���Vm�p7io����Sυ�����n���O�Ƅ�ܗ�k\e/�B*�������#����~�쯕F���դ�����XY��t��Q�Z�'*�R!~��VX�L������廨�_���x {�?Yl��`���T�hf�h�,�}��� p����a��ի�a�+�-x�.��c�v��{+�|���ķ�/��-)�D��������W�����kn�\Bc5�$�qpC��;��`��'1:���{��*4�59;�"_���p���k ��(.�עT�Q�j��?cr������ǞΝ6���պ_P�M;�n$�	��c3ҕ>�rm�mǊ�lO*���P�{`OԱ��Џ;���E��-�_��J��@�����O�lg��+\��/W��݄L�"��G�� 1�Y����@��^�m2��k�ӎ�~��.4�S0�(D���k��N>��g�!�3�v׳��̟+C.^v� :�}]^��`�Īg`�7�7�}GĂ����8�ȗ=�4�S��zBف�ʰ=�Zt�}#�>�G�nzR�|Y���#��O��p�y�%�o��1�D�ʭ,��Ο��.dϯ���A��J��? ���jb��͙ځ� d��d��?kk:\]�r�Y�27����Qㆪ2�<d��#l�M����r��?3L�h�:�ó�k" ���Bn��;��PFW��MĠ})#�~�O2�~:ˀ@����I@�MAbc�n�.lGD۷V�/������Ĥ��������v-8Wv��3z ɞԇ����JS�CK�l�WIOR��'���K�+��'�Ov'���5�$���1�w- !BM���j����\)S�Z�Ȣ�i���I
���}�D���$d��z��(�w�)T��"�֍H1��$������T�]�������c�^L�R.�oJO��2�����C�:��G�"!��P�Y	  >v'r8�EͲ�\8��8ύ��������I�$Ķ�%�$d8�չYc���������, �>b#�t���O �-��{���ŁU�s�(U���Ar����ؾ7u��J�/d�y5�.����ɻI�(Y.���p��}dB�T���^J#@�v�Y"�2�A����dr�����:N��~�}}+�7՗���W~<m,�暨`��sm��e���seM#��k҄t�{���⭉�^�&�¢�wy3�\����$���9J�C{�YWL��w�5.�����v�x�N��&�s�?h�|;�Ʉ�Y�8E~7�F(Y�:f�=d��
xx�.��g۵�c�~�oM��}k=X�b� hw��q�.���"�	�Q�}ۆ/����}(Vc{�ʌ+O�v!�T�D��K[~��������9Z�
�j��\pe�σ»�� 	��zF��}��}�K�O�� ބ �;^�� �ʚ��˜ƅ7,~������i�{��T�B��!%Hi��<����#D/*���L��"5�8�m��|�	Ěe0kk�s��� jU"�o8|Sݤ+��l���/S��^��TIOU�I�1#BE@g3;»�%�gj�z3�<*��}2!E^b��i��W�Z~��A�L	`���[�%=�E�Z�&���NpR���wr�/��&i݇�A}Ds�=w�Ճ�����K1�����$U:<�F�C���ZR?�q߹D�`4!!�O$��%
����K�.�Ƃ��1��I@�OU4\z���Y�ZE�i(.�͘��zr�z~�ə�����|{'v�]>����@'_�}�v�n�O�y�|��G1K�����i���1J� �\���FBc�@H��v6n�6�_�$��|M�Z�}�g%&�ܓ�T��ø� .s�y9��p�_��N�A��`NS	L��Ep��;��������$�|�(�G��a�-� ��:��?����$�������Uy{�T�4����]#���B����ou�+z'��h�2�G%����{��r��
��3���� ׮��pi�p��9��ei�����'̛j6�x^�B�A�E�F�;U�L���c����־�P�v�T��(J�Vo�F0Ni"}�		��%��4J�uy�]ד��{[��N�N���"�֡�%��G�v��(�aN��lSy�WP�S�Ykab�_��E��f��t�DCx���/|�UΖnl??���?�C>�4�*$��R�畬����O>g����B�����$�g݂��7_X5t�=ir���2I5��y�u��^ϕfv�5��s��&ӭe�F|�us��9�YLJ�lj*��_�6���?�W�F�r��`m��Zf�r{��Q�����9�R��|��� e؏��n,�8�Dl��w��I> <��C�(޸f��y΁��*P�ƑۮRvf}{��ߙa��D �l��Z�� ��F��O��>5	9u�Ŧ�%��y*n�H�dؠ�Xo?�?�Sy�,$���dL�T���<�J9��L�m�Ķ�ȑѻ��_���&�Q�֡��}�k^�C�U��ǳ[~��9�i����2���{�y�]v�Cߖ���2�_�2x�Ӡ�Uek3����lE�d/6:(���	��D>aˇ��?U�QOg�U����Z�`�__�����D8���j��z@%$L1j��R0�������D�I>:o�o�� ��
����bO�J~GZ՜�g*��o"8ɋ�#oX����hԩ�[� ����y'a��Bǹ>C;���o?R��`]�~��\v���B�t�NP�Fmj����Ţ��veY�X�\�mO�i.�xH@��$*j�U��@�Ee���V�^m2!�8k��hY�X�k� M]�j�2ɍ�9����O�i.���z�Ĩ�,�a��c��L�#��aϫ�qk|�4�5��*r��a�s$k���RU�-Bi��­��2�����sG�줯�·򠝶C�=]p=z�d���n�Ɛ�7���L:�х�+���	��5��A���]��W��Y�6�>m�3�Y7�P��?f �ZF�z��#����q:����j�5��X}�Cg�E���˙/�������V��f.Ԭ���	�]T���=�����'��QaNULE��r���i�Ӯ��NCt�ECBF�$Ļ'}�>���c=�硠��DI;�$RR�ؼ3 8J�	�%6-D��RʀTDV�*�C����9����o]>�%J9c�.0H�cU-�LHg��X���બQiv�*����ny�|�(��+�f�Ϸ��x��ɸ�������s��$�L�g�)�@Ͳ�߱JA������7��졦&y�wU����^F�?9<Kȗ{WA���CT�9�I�ķ4zyba�l���{�g�U@q�,ۮϭ	�"qsO���j�<~B|��H�9E�ةs|;�D������AsFCH n���m��pS�^�N\r���3(�xg�9=�/D�j>CyK0�R�ܬ�s˿0�τ�b�gƂC%�R�}�!T���Q^�b�iD�B�T�&���P�/ђ�'O�b�����r<��0�AR*,N����M���Y�&��W�Y~ӟ�kC�i��ovDg��M.�v����!�g�LR������f��x��.�p�4��4����$ZU4�#Lk>�+f��{2�j��o��ܥ���`2Ы.��^-�ni*Q�2�vR57?��Z�lz�0a�(���X��8Q������qnӮ��ª����gʺ���M~!���o-�%������{P���Z�iӤ�_�����V�/�!�Rs�z��q��W��l��r/:�v�z��mp�V�I�t�ɓ���ӷKw��p��A+8:d�.qc�<9��%�.����#�%�C�5�]��A�Q쎍Q ����l���҅��8�u8�AI��d���ɟUy/���y�%��O`f��E#�d]	��O+��?{�#\��C��a��d�AP�:+��2���&y��sqr ~�ZP
8�j5��B�����%�b#�V^��ڹ�ʽ`����z�Y��E^T&���!<Qu���fU������GZ:��q����3U:�+�r��xx6`��]`&��K�<�L#$��)ו�V�5�A�F�yR�\�Mj��3��)�u�	�����}�enB䫁@Q���O������aq�%�����_�otN�]��.�W�	7<�:e��\=T��M�a#��86hq����)�˩,���A���fU(d�d��x|?��RC�XI�{-b�� �7J�1͝L��)��y�z=;�@�t��h�Q�������(<��=7����{��A�3��ݫ���?� �1q�\�@�b6e�o��rg��x��������G$�h�VJ�_�8B����{�F 2������Zzկ�����9=�^iR�;�`.�Y�X�S��ɠMo��c*�G��d��mE�d<�_<�����L븃X	:,�b~c9�>l��X���;�#��U����${V�������U,�f����@��] ���d��Be���Ԡ	��<��S�$r�$։�Ԡ�i�L��dc���i����g��_��~��wz��x���MZ��(�X�o������Q�ܻRN%�s�x<�U)),k��n��S͹��3Ʀ5��z�����ʣ�+J�����Ú)����t$�8�gu� G�0���WX��eG��u���j�S�Fl�����+�Y<����3fZ-����b4��d�AɁ�����!�o�<\	Ш�̢8 YP����C��t���$1ҋ����]�zkF����\n��̀B�ֆO��\T�O�oL�S����tv���1�� h�y�^�0��v��!#����ț�e82\�
+�!�UQ�C��8m~�eaYxZ��m@��U6%!i���.�`����)�D����~B��"R��'�h�ɿٲ��U�Zmr�p�]��~zz��{ (�3;�n>y�7��;FxN6�@Pq�?�6�/t��ҋw��h�e=��2���>�ڈ�zz����ëp�"�g��*6P��2�^9xe�3l���� �<y����>+�I�ħl�8�2�z��[�����V���P�w.0�������cX;J+���?�l =!��`�L������z��Z�-JWQ��P��Џ���}�M
���[�.�-L�-���I�&c��.����_��%�sy�"�DP�X�j�?,@�Us+M�Y]wǧ=����.�vW�9?��Ok< Sgb�6���'Z� �þ���6m6��h	�^Te�[
5�g�>��_gx�:�Vn��WŊ����1G�L�u��H��--��2���eJg�RB��`Q�6h
���)������SS�x�bx.r���6*~��M��}?\�b�8'\�0��r9	��=���<���(<��381�e��?�ֶ��۱.DN=;m�l4;;���x���O �������dʪ�������=����9j��V@��l�����O�M�[�Ş�xRj8Y~���ra�������ʃ�-9&�6�.�I1���&D�4�����?�Q"?��L�4vN��8ar����$x�F�&�H�"��_f~�Цeb˼��f��Cز��BV��G�v�U�������NJ���8��r���F�_��R�]=����; �5���tG !���/jp��q��nK�TG�Qa���?/6B|���`Z��?�����%�m�O�=8�r�?B������}��,���m�VwXׁR�'/Q#i����i�i��+���p����RBq��D�o��)�n"���p:
B�v��BLv��o�����s^X^��c�,D!x�:�	�9&Ĕ���v+j��)�-g-]r�*
)XtHvl��OK��Z�!s3�V���g�����Y��kתk6J%?yn_����l�މ؇��+	�-8��K��g쬫�
�d�����c�@�N<rY����=cs;�1M�7�L�aдl���ȅ�#�(o���1�������w��l�t�D������rޟ��ÞǬ���&#��˽��sN�R <��:�W�E�s����s�i��S� ����>s��K@�K��1&)6�`"�ڌߙޠ��,/�1-� ~s4(P�qgʊ���ݗ''U{ƃ�>{Wl�� �̪kwd�[����1��8ֆL�hM]��E�*����S���E�SJ��<�2����q ��#r$
'�Qs��t���t�{���,t4J�|5EX" ����(��hK��!Gz��g���ӣ�����I�&�`I�zqQXj30ZKJ[ui\6�c�[�%;��+:��o��?�*oUS3����@,�z���'�EgՏMx�QĴcˈZ?ݑ�{˘+���>���qd�?�qr�8��*[�j�!h" A���yE��V�P[[լ&�ß`Ftvu.��'F{^�d�������M���f�I=�R��z��zy'�����F������p#aA�7��l��gi-�>*�
^��##���e}�D���<z�3wa�Y�r��1T��#�n�����ߩT�����͟���ú��0�F�����m��OܦӞ�и4��$�B��_��Yo֯�S����P�{���L���9i�Q��	v�S�6=жkP��=�Aiq��w���){����Dk�n�~X������������
rzfi�ՏN���*2tj�P�6�u��|eo`#�Ǣ�#�-�O�+�A���T�=�^�d����{G]Кa����uS�:�=��I�a���hӻ��F��3��]{6��n�Xe ��'~����7p��$�Q,��<�nl�� B�铻仆h���֓��9���~gj���F�jŠ�[}	��#,��~w���|v��l,���V�+	�LQ��XEl�aC��zٚ^�y��~��E��~�ԗtBT1 �z�*�Yc4Gl�o�?g����B;��zH�ұ����H������H��eP��C� ��jy�4��/I���
&����l,P���Nj.�u�,^6BU%�ː!�(W>[�>6��'���Gf�G&1K���Q�+��j C3׋H��wC�:r���5�\a�	EHi�$�(E�s��e�G*�It,8`P�%f:`0x	l拰�k�m(��T��Q&��\(���nL�8O۬��\ad�<�o1���8t��3y �7D�z�B>�!sLE}a�(��3�$�Ds�]6�M)�et�d���D1T�_oʑ��^�=}8�uL<�����d��P����h�7/�qD�|f�Gsߛ�����頃AA�xc�,0\��������y������a������36P7k�;�?[��*��=��7��W����r��� �̮�O����e�3���=������:m\0�H�e�	{��_Q��?7R�z8"C���.�J'sP%ǐ��ӏ�9�P�\���+���(�z_�ΆQۋ9ұ9s�r4����KJ�°�2)�cyM�T7&�u�w�<Q�޷�F?	ݫ3K�lӝ`�5R���./|���>Ԧg:�;ȇ��������"lm0f,��8K߇-��=�|A��լ7r\��I89�H��p��-�6��4�l̢51�7��Z[zo��� H�܏Oo�5���\�ȶ���!T���e�Y���j���g��R��Oе��j�j.�%�U]bP] �5���!Q�h�8�-�jwg:s��P P�]_ˍv��K���>���`����$���3��_���{_�R�6�C���sH���JqӍ��m�7 $�m/�l.qs홧{ �8���MF�CU�3{�a�S.HŪR@��&
���wiI󈞾��1���]��a�W��G���S� �et�YBa��{�~�,ܮ-�lO�ld�G���|���h��� ��n�? *X�{rp#��d��MB�@':F��]�̚w�d�BZ\]��E_[�����vC�����(`�V� u�̱��7ط�v��s�8�7/K�oMi�i�wq1�$3�Μ�� �q�y�7x�u�D>PC��_�_�`i6O��̷697��K��"7�
 ��m-�&�M�'�Du/��1?<�D`��h�����t�!S�2��r%a [�x��&�� p�N]�ezYGPR�Wg�%4i;�u�����C[G�������).����:yY�������; ��q����nk��ӹ�E	�#�
��u����?:��HaOn��t�]h��Vj��Y���7�K�t|��b;\40�$n������zԶ��w�KF��#k N�yʙ�������Md6�.����$������!��3���L�}�����~Z1�;?7).M�L][��Gߨt:w�23���<d4�;a2��������^��'�|�ڲh��x:��x>@�*aT3���Z�B���"�Q��GjЪ�����'_�����RL,�%��I���R�EW�H���-vcV��g�dc��1 �M�M��<Td�S���(�)��hQ�~0.��6z��&�b\(r_|�R�@���&�\@wH9�H�!'��\SI ���G��V��9��iumQ6����A1��'&)T��LγNM_��%�v֝ˡՈ-5�.��zԡ~,��GV
(KJ���|������ ��;�س�as���[���ؔ5��>='���g�UG��� e�G{�ژ:� 2����	M�q������IR��i��o�<rd����ŏ�b^T�'��Av��8H�'$$���1�� ��"`��n�1^����a�l�7�Q�ͷ�M��5�>�6m�װ��S˄����Yꊪ�G,�� j�����L!���(ݩq?F�*�6^Gx�#�Z�V/�p��g���@YKV�A	iP	�y�Ӹ���zIR�}���t/��C�N B���'Hx��&2�uZ��L�� w��љ������/���z�.̆w"׬���R`��73���T�4_�9I���������h�E����k,�SI+�<u?N�f��*�L}.FZJ++�~v��)!�K�t���U���Dr%��9w�s�?E<�(ѱ���|�g����pj�Qf�8D2G�c�M��|�;�E��?EiK1vBS�oD �~"O\ v�>=�Vֹ�����<}'��d�<@���2Ϸ7�ʡy3��ZS�p)��pi̱�g���PFFLb�k�j�[�c	M��ڽ��ku��c��wP�o�B�K�Z��(���9��ۓ],�{�+�Ԋ8��CZ���K�B�"}��L�>_n�|
��[%��[Ms,k�}��ɋ�;?�0=:L�$f�H�39_����qH�|�e/�``D#�a�(�)x_ܸ�d��M��vT(�#��(]�j���+>�qs��J�r���HX�Х�7�e�3��B�dH�$��{�J(W�*
�凇�];r�8h����] L�|�߄7~��YYΌZ�L<�N.�2�	�3"��)�G �P�ĵI
ѥ�����/�׫Xw}П��q�}E�w6��PR��SW���w�'}Y-�!'��� �i���Ж;�Rki�C���j���~%�y|�ibjA:�Bk��D�h&m	g�	F��� ô�*,?�{��!xt~���W����y��`��.��q�:�>1+������l��C]H��wm'�h�w8�&��vN'<�P� Y�w��i~�d�|� ���՜��#MW�X��D�h�� N3����EU���>�׫�)I4��L��ᴹ(&�4�2�,��쁋��y���X��]/�@�����N#r��ݰ{���Y��HGP�WW1;�ۊ K��@�r��M����z���"zE�!&n�g���(���h�����罍1sz�/�Ϝ�l���Mz�9�Կ���	���S'����k(�gڊj�k��w��Kj<vd+�/��i��hAE]�^�떣�'G G�գy��J�܂Bm@:��)��S|�{]��w:��N�k7s��)���J��Q	<󚼝ëIR>�T��Hf���^g�����]��߱1`$tEc�0�.pG?B������r���N��ij~Y�56ӻ������ђ����'<�Χ�]�)o�c��`7�s����uꇉ�-�d*t�@�t�4�jVnx7lK�Ĳ���I,0�w�̑�M����֤Z��,�.��>�9y�tmcPt�>���7YyRO�43��
c����Z��|�!��}='_W�~��%kI��	��3s{À<��o�!@÷k��g3v�(�l #��3I2����,�r��A���n�6S{���|iqڵ�F��۔�^땂�b�/��ɭ?'�����&1�"'�M�)-�*K�j(g�DG*�؉P����-h�l���h�\��VBWd��TM�j!7�4�G�l�P�2��S�e�J:@X���5a�-���O(vf�⫵��H>�]�=Z�)vV�g9#�K�<O��kU2O��D��:|�y[�U��1�K��r� F71˦��W=���ʘ�T*��o�U9�r���v�x, 	��U	۟����fG��� !ސ��Pt$��޾/ݺˑ�s�n�G�����x��'Հ��/�+X{���yo��Ɔ�ÇvD�n���U4���t�_\k$��[yD�A�����������S>�Nd��P��c��YK_g\�P�1j�(P��nuJ��EU2��Q#��޺�/O���iZ����-�rq+�s�|t����-�|����2g4��r_m�wA6�D֭����q�_�v���~)'��{W{���ܨ�3�ֲ�&}��k�_����7QH+<���i��: ��NO��x�^��_M=�x=Q��[�
�V�w�Z\�}�`����jө8��I+�Rh����H��ӻ�8o��z��$8V�VT�(E �*��a��%f��J��XNB�U��9a���)�6��`}����@���S�O���U�,��"������ ��񖨔�iI�Ӎ>��OĪ��mk7.���7��xB�N��n�jOIQ���sh�Ls�&�-�X���2�ث��j��Ӌ���_�ٽn��,�*��H�#�H�K���S�Ým�D�@ژ��~yi�/�p������� �)O��z� ������cb�<%�B3s�c�ޟc�:��b`���I�}����%,�!n�!|C�c:�=mdO�5{K�Nbz�b�;�C烷�e�P��d�mԀ�g�А���#���&�'�z���;p���ū��E��ĳf�z	fm�g�v�g	
�{#r<^��9������M�%�c\�j˿<�]�=$�U8Y�hn��-&�[��wJ�C�/�g ��P"���n�7//���P�;;��8��*?�]�e��V7�T耧[9-hjR���*����u����C��HGg?&�n�d_u2 �3�_�g�4-0.^L�]�S�tX��,¿�S�{1�l�q�.�ag\�ˤ�Ŗ�E�ՠ��~�����;q�cV� ~�O"�@r��0����6�?`Y��F
��5�E�f���W�#c�����^�y20Mf{
�����.y<���]ʒ[�½�J3�b�K�Ӄ�H)��n�9��kqX��������ߒ�E�nZa�+����6+{���t�6�eQ�eǥ���uՍ��}�ssp�D	��"x�ϺD�#���hl�����%����%t?��U��c�4Z�\���Wd|I=6~+C>�c��_��.�����1I���Oh��g7��09�Q�#�-�&V��Q�F��P7��.i�"���;��=�RF��x�]�қ}`.r�,����r�0届�tP�m�6�#����Aś;�L���ac�Y��WVMw�x��R�3�Y�Tb�m��=S@��4rݚ��3 E�I����/=d$��W��T68�fo�!!0���O�6����l�1��֝�A���{�]�:Av��e��C �c���O�=&6 L��T�Ƌ��.آ��Zr��y�� a��=�ƥ磩�X,�7ݻ�V8"���k�[m�_���v�#{�N>�^��j�S�����p�n�6!<��.�bp�j��N�t��u=����O�����߷���hBa��P���{J�e�b����h�S�QZ��	��u�{��^�:�hh�:d��P���R�1�p&��g�>WL�j�u�;qO����Yy�j]�|�˻ij^�z�QksX�z	R�~2�J1 ���� |H�how4�c|��(�O��b����3���-,��a�K6/��^�V�%\���2/@T`/Ŕ��
�B0�jo�(�d�������" �"" ��uQ
�n �_���sTO���e&s�I��C.*$�e�^>H�'(\��/�0U�,���k��G�i̐z5Y���䘃~ǩUo������{�F�L�1J�J�2� �R0i�2�h��S�ad�`�-�����oP�Z�$�d���A�&qh-xl �g'�AC��1��8���W�|���5�+u�x�R��m�#�C�$��>pQ����KJubg#ȿK�7|�}Ŧ7��G���KV��y��k���
�fUT����otү��@� 1�l���������f�l��@4e{ �-7����=��*������6~b�>�5�S�1���5���ek��8~��#a+ݍiE�?�R���h��/fM	C�n�Q!��G��4������w�����+��px��`o��Z�J��y�L�>�ul�RA�h�Z���W�s.3s�_lcǵĀ����I"�Zt+��- �}m��u�6^ޮ�����[{?��My�Vl�*�1��M�S������揿μ�D珗j�".��و�_o/Yk�|���}w
�F�P2���&���V�`��*�[҂B�"2�Ʃ1����8:MOuL[׉�$�XBwvd�+�^�
���Z�+��N�lOn�!3�.�̾8�J�20mV��\cS��<�T�ZN�La���m�U�
a�E:�^e��v�W���^~�c;��s��o+W��&�[]DD����*$�:�ä%�/M���Ev6
5� � ���eF��� Ax�@|IDF ��Y�tN�(3��%a�]�����v���8����a�� �fF��"��ڪ�9�3���� Fj4�E�������x$!�0���(Җ�|�wI��T=t�^9|L c��"�--��)[�/�=��OG������9C`*DPoI�3������Z`��I��p�t'���p"�������_!>):�%Ibf���xY$;AH�1-2�$T@�{���Ta�|��iav���l��I�!���a�9���"*�R�.�G���%3�e���µ�a�2���f�D ��A!S��vŵ'�����[�o�݇13ꉦ�$��11���c��H������L%��g[_;�:W���{����<�t��bn\b� �urz�z���P�K�!��⁺���������;�x��XPDg�H���!����!���*�u�IAsg9��W7�S��zZ+C�#!����0��}Iݸ������[?�&��rVA��t����Y0:��-�ќ=�[�X��Y h u�pγ�.�_>YI�O�ܙԢp�b=�X&���|$|LZx
��SP��.ӫ[}�ky��YM������1�U��ec���(�6U�[r#�/a2��ԟY�x~��PWر/��[�ض��y�5�ܚO1������0l��Aҥ��.L�j|q(�v�ӌ�[��vo$A��/�I�8����c^n˟3�v��ğg�� ܢ3 O)]�1��Wa�[�a�'<�5YD�C!F7��^ӂg ����E���7����q����Y@�T����[�-)S�H�fe����5W՜�/�@��=�Η��e�H|�&B�'f�l���S�y��@z���w�z�[ִ5�
���<�3�/K����z��`*������@:�'D9�<)��Z��v��~4���3�".@��+2_��$���ᢪ�������;��������=ù����u�#�RO#TEAK.u|ش��#�mɐ�Z����i��&���ab#��=�4 ��P\za2�'�����;���7��aT�KB}t�pr�w�[ <�VE��$�hR�_.�?s�/��#��=��Y�k��8������}�"��:�&��|�j�|��,Bb����4I/do��U��H�Jb����_EB8�?M�%D�Z�/VB�Lb��\��mx�Y��5���«O�?:��#����j��BdљPئ�-�ss ${i��-�eb���0җ3���MSd�c��6\�����j���`k��Z��l$��,�w��tԤN�*��m��ap��>WR��2�%ܖ���;�X���023�-�ؿ�ʄ��#�1�o��OD��\��2��qc���Yblʪ}c���M�f�b���Ʊf�VS4D+�U��?�/�H(�������t}����*t��_�B�lպ�LS��x&:���`?��u�e����WF6�-���JZ`Gq���!Td\��Q�͞V~n�w{V�d�8��=@���S���6��*UQ��L_@3�M���AJ*�w��H�~�����Nm�4���Ț��#2OUڝP��zJ�{�Djg*�cvO_-�(�0���U��0}XS���ўׁJ�� h`ʫi�!��/~(�l�t�8]V��u�CX�W~��xs%���AtsW9��qKzm���Vܿ�Q۵��0m��ڈ9�"�B{��m
\�2�Lq��ɖq�����X�����*�4�ᖇ����V2�ϋ�� `�X�*�͟�.r`��W%U"(�N�a c���ew����";���J�i[�)KR�%�ј]��tJDf/7j��S����MN�����:����lˣ0R<�o�n�+'Ӧ;9�s�AT�+�^ҋe��ʒ:�����E�)|�|�Ff�Dj���<aO�`���M�,���m�rK,�E��^rY��?�R�&��jĳ|UID*N�v���<�����wY<�3А��t�t_���In��l��Wš��2�'�[w��p=+?=�˨�E�W��E7��\�aZ&�{��FtPq��_�=oĢS�Hp�l'{���B��l���͸�Tf�7�3g^R�,�~�X�&w� W��������]�=�{�jG`S.�d}��oˠD����x������I����#��^PQ-!�S}�;)�,`>��`E�a�����L���G)!�g7{��.�CkY;������@p�~!��t�?�j1�8��G{�j]��0��
���uI��R����=�����]w@F��{`""���S�"+0x����
�I-2�r4�_I�
A��/��F�AO��nÐ��|&��m�
2WP3M���D��bA֞�Ps�l�a^���7M�h�Ff�T�X��H!C�v1̡���ن����6*�y?P���Tr��e�^��$�
6�Y�B�Z�Ap���� i�����7�j�o�w9�t��{�.�~z�r�`����X�&d�^۽�Z�jHI�;��H8m�/�����iI�;C�yϬ�VLqWQ�Ϲ�~춊C�Lk�y���W�g��U#��rZ���c�5&�6��庳ԏ{-7H&�����;��Mg���{1([��	G�YSF39��_Aܑ�99����=�1�<�ʤ��E�/���h�(��z����KrS�N	�v��9�麵�BF@�kp>��� �z����s��{Ď�&l��S���9�oϓ�8�}9�9x��Pdʦ�∡87�Y6VGl1O��k�/��L�ʮ��k����?.��I�����^�J7�
��l�ܛ1�*'�LȪ��I�Ҧ�J�Y60j?߮8�<79�ˉ}���NX�"0@Dr�l�!0�����W'��J��$a��lc sٱs^��Ӯ�=#A�pM	�����҄v*#w�!�0���d����َH݅E�zE����]��@4������l��Y��x�E~)�[=X��;[>�:���@BK"��%�|�Y(/#,]]���Q��$J�Z�#ז�tPx�r���������`#�xף��=2��������h9�J���r(.�:� �b%"���Y�[y�C��Ⱥ-!ej��T3bZ�[N`��۟D�:�5Y��]v�)!�n���b�^�H6\�#r.>�`R>|�{f������c[@�{�]��Љ�8�D��G�Չ�&��K�.�j��i��'�v�4�M��a73Apw��C�M�ڍ6���+k.骱��K��nK{׷-��!�ĴH8gbH�.�v!寖Ph�- ������b	'�,� p���x���E��ra��2���bC=�@����FՐo6����|%�-��>���-	���˨)CIgה�q�)?^�&��{υjF��? C�,h�D׍ĵ?.�x��%ǥ=1�w�\I�,����F���s�F�7��&����$�i��"R�wp�}*x'��}�PU�Z�8��)p?kq/��;�l�z)D"��.��aaz�-�aV�����a�
���AeE��oE֧����t��-�酱�_'lrb%����������Uvk�=1�x�|�o}�h=1��80�{{��$��^Z��һ�S�l� ����\Y��R@#�ѻC���/<!IQ�9��4�P٩��Y]���.Zل�RI�ڸx2�l��Nv���e�]�]�������\4��v"����k���'�\橳{tB����$�P+�i2y �	��E���"�KbZ��}�~�Ţ2��|��-���C|.�<z���E��vK����y�;Y���zcz��4��J�㒯;����R�`KJ_�rŁxۈ�{��wi�ٴ��}Æ��^j����B�	�2~�A'^�$�.x����,�i;$�i�����a�&�V�\������O=ß+�47]��t�tVV I�i��	��湏�z����f�6ޤ�&��/�|�Qq�Iц�u=p�	�\�w�/�35'�×D'�h�Qg�M�t�h���ev|�Iu J�R1YghA��ޔ���eF�y_�N?`Zº;D;��<dg��v*�HxΗ*Z"6i���s,�L0�S�XB�M����;�1s�'],(���F�4<�`�sӼ�D!8F��\
r�C����ʩ�(��)�Ի��l���l�vV�f��U�B
�C����U�و�;�!*c�tY�h�7�����A3CgOI�,`v�rz��|�V�K�p�ĳC#�[Г��x�T��b�3�*�>�3	���Ճ�x�ۀA��9�pYw�q�S?�S2��8�5��#��� ���߸���L2�����R�[)�ha�I:�!'� S:[6G�k���z���>��;�X�R�+Q�5B�+���W���#�����T�W�P3B2��ݨ��,�~�@X�ŽR����.�4GA
z<D�z��?= e��&�w|Vq���G|h0�'��e��M�4�@N�x@���xh�f���M5	�&�h(i��ŷ�7(��������x��֘^�X�ѐ+�♬��a��
SS�f�Lա��g��\Cw0�SU��A:ut�k[�0 �YKB�e����d3dR+�>c[���0oH�@0v5�C����V�F����e	�P&|��o~̓�`��=���W߳�ZpF�/�k�6"��{�.D��T�s��n�د�� Ϸ�H��'N�D�vn���_��;RB���8ݱ@��v-f_�n��+g�g����3��u���ۆ@ETP���3xT��7�`��pt�g#���/�çиD�t���ɦ�Ƨ�2�����z
솾G���	�lR��z��b0���C� B[�y�_��@�hnKݦꕶ�GfW��{�Dk�v�߹%,+���-�ﮁN�<ʬ���=����!�/�P�E��[���
Q�OڼFz�;���-լ'6�am�����9�
�!_Ԏ�����	�Q�oq��\���nLU�RnR��Y>��#TD��hl>��Ҋ�P�#�-�\�[:���`�	c�m������)+�����J��
����O#�Ó�<dt��5E}����Aѓ=��c���❣�~��~�]r�0l�����.�����v�#Q<[	�����)h�pH���f�
d:w6�~�S���������n�Q�������kP)�i���k�	�L��������1�3I�c�����-j^�~=�g| _�`���z3� [�@%�RXy�=5Ђ�����(��}n	�f��eq�\�Uz�n����֤!2Wr�F�.>�O�F�LI�����}c��Y.�b���$���j]�A�4�5}p^dt��^ C\B_]�E �����9�i�69��6��V�)n����w9��&��g\5����A$��ö��mZ�\^���|���6,��z�p�ӷ���΋�@A�G��[�s,�����T��_n�E�쿻h�Dz�����"0� Z 6>���2w�J-3��]�a�=�aЈ���q�+�ö�~V����hn�@�
-��ȟlC�B�\��At�l��m}��]�S�|wǣ�f	�̿e�nn� �X�uBW�bng�Wl�	�1�R`X�U���·����d[�t���b�&��3��eQ �ƭ��?,Q Ԍ��ȵ,#x�����6=�;��cw7�tl@��sŅ�@�+�R��qFd�k�/5P�{�'�t���D�!�ς��Ks%h�%k��m��M�����d����������l��>�b�a&�� M���\Rd"�P�$/y.��t!Ls0�nn��+J�_
����:��r1p�_�1E�F%�!k�4}���ŉ[6o�iN��j���~�h� ݝuҴYn\ퟔ0��:�F
@��>3��m�qP/�Q��緦���)JR~8���N��+���^`��)���_b�hY�)x��X.�L4	P���q����X;����K�i6q�,�&�w?�����!J}�H�k|�����Z���؄����_`5Y���q�Y&�A�@]Rհ�{��FܷiOJ B9��؂T���*�|_��<L�*� ����Ҩ׈6�~��"%.�<����>ԅ�4�4_u0@0��%b�����g^@�8���f�����v���3ۙ��
<�]�E�����F��k�h0�HQ[4�ך���e�V�|V%��I�x�����q��7:�ʼ)؞IO�?��h�#o�v�q�؈�0�q���E�����θx�d�{�`�(��������YS�I:/K�t���������-$g\H4 @��������G�YfϏ���ק%�L�)r��=[|���������)�V;uи�� Ckf���&R���c
T�#��j������dL�/�n��d�pۜ�&d����n�m����Tl���� ޖ#@c�*n#��i�{��ϝW��ING.�n
&�p^�/�er�G>��(�*��6�JF�O��kkIr>��$z����3$	v8⥭.P�IN�O���]�@�����������f}�V'��K2�̬-�ӫQ��3�ʼ�]���Z+��Ej�H��ot}x�O}�y�E�p��Z6]�C
4��K���F�  �2�	�J�I9=��P`$|ߕnk��ݚ#reS���-<i��g���5�R!ö
0�Է;<B���0���ѽ	_�q��_x[��U*1O�'3$��-4��E���7˷�=�p;��j�m)�,5��8����h�݌x2-IdA"� O�L
�s�+�@��q�5�G���U{�;C���/�:��	��[��k�龎�b~;�� Y�x �� B��T��M�dm�2 1�y�����A-)I�z����w����y��c��@|l�Y����z�������㽮
���TUn;�h'3�G
؞t�n[�Z|Aa\���[�'�l�������(YoL��	�'�ƫ�ӰkCE����Մf��n�馮h�G�+���C�+�-F��E9�}�ގ̵�6�6:�f�CK��2p��J�;���Q�&A�������#%��(�ĺRub�&X��c�Kz)�31b�҅�ǩ�hA%AS+�Ҟ�8,R��ME4�U����4D�P�\���I���k:5/�.��>��e�_����Uw��aDN�H�]�+廃��%m�V��� [��ioŲ�eNf��b�&�vy�q���&#��ܖ+�������0t���|�ߎb��Ob*WI>��R�U�T_�j�ֱXQ<\�*�EH���Z� �[����Hn����<��Qꢄ��˷�h7�Xy*!�b]xPpA*�	)�qiѺ�s`L����3E���f �ގ�1��⧿��R��hj�?�޽4Qm=���CY���%�X�H�D���_�%5߉,zjwZ7��rrC�ףV꒧�J�����o������}����L*�~J`�}�����Q��
t����?Z�=|�kc���mX�~�`_1��[vG�q����Z��e^�4��K�*VO�q�QZS`v�q�l_��������IГj`��8�Jf����M?cf��C5�����Jg�������hcFd�7��L���9u2�j:n�����Pky��{���5�p��O�o,P�Q/�T&�Zi�a*e�u'.�a<�ʉ)#�/����!p���#��`����x;��_¼���^�r��m��l]\�8����U˟#��F���{�`��;>��Z�\�걊�A�̕���Ym�t���I(q��_Ct��L��Ԉ�2�xQHV������Q��H��@�������	rv�p���W��m���E���=��P�ǂ~梆�J
�pW�u~)W��E�CqV���#�<�+d���Mk$p��ž`����}9ǘV�Q��y/Lk�5.����v�>������0�]λ"ׅ�1X���b�(�����c�$,���8�mYQ�J6ٛ1��y`�m�yGJ�"�}�m��Eh�|�D���IhU!��Tp+-J%V���a���$�)2J�1_�����q֛�]���Sz��N��=�s��EI�5�[1�H��r-�>N3˗.�Dq�D^�*�c�J�6�/�;���P11�S�?j�@>^�X�*4��9����5�Z��ǲ�m��<ɿz�xH҄��{���֐���)��H�~��W�ʈ�\4�Ԁq�#V%��:��]2����r}�D���v��6��	��F�[ʋ��4�!bK�?���(�x��U]�h��Uǣ ��]G��:�U;�.����F��'�ʘ�.L��	�zB�,��p͞)��H�+[�g��>�Ɛ(�i���`�h�	vG�h���*�>e����_�3]U�i���_nF��#{�T�w[�+��T1�2���8^����:!����{���b�)�cP���_�i]#�
���PoJ�0 �f���0����Ѩ��R����`��N+'Q���n�H�p+�b���) c~���{��i��I%�����_ǳ�B�<�ｉӠ�����I+�9?����G��;�o4��vy!=OzZ�i$�"����Xa�y�3���-��.b���tQD���'¢��4��d�N��f�9*�<�4�o���</:��I������7Y�(H�+A�1�s?�j��W<c��q&U�WQ�H
�F����
ւ�+|�JAݤ�n�P���?�����00���%]�a5m]�7+�%�zP�7S�6���w���I·r�*�\2�g��teT-f�]<�\"��+�[Gk59��S��1���se�Ă�Ř2����۔��ď��O��U���^DL>p|�k�.1e�4��v�p�?�d�j-�=�F���\xZ���K��烺h�m��<�/�'OsW^-���o|IC�R瘘X�K3��12�U٢�p��,��J=�*[zDDy8#1�r�|��2���Χ�V��6@�EX�w"��_݆�u��4��G�KMd~T�^��CYK� ��8c�׏����_��WG�;���� �O�h��-�aQ�}��L��b�Ub<�'s�9�"�?��B��v台A��*�c*��I)-�w�#iqE�y\���g����]�P
SGǡ�>��žtĮƙ��x-�s24�Y����G��1�.�m����[	K������"�F�q`=.���	;f�T�O��:��`7_��V
P�ܾ��~�m(��P�ormIC#���Y̎������ߛwW��es-W���o�^�,g-h�P��#�����C��Ɗ���R|-�KdQu�H�.VU��	��Lަ	n�^�a��c���ִ�R�1�k��iR\��ć	�����Z�����T���\�M
�RߦSh�jk�.-żk�O���vP�@�e�3>����Ӌ�\h ޱ7I����N��C�o'
3��������#&0g������3�B��)�g�ϓP�� v�!܎�N��z�������0cS�|�|�;}���n��c+/��XQP>-P�PM{;�#�}�����̈́�K�+�����B�2���c�kYlg��o��HÍ�I�*���}��?8�_ʓ��򖉴�g�A~�c&a'�G�g� ȁ��%�^���l�¯#'�FF�>�J�ҳ�G�iT�Ch�-��Q҃>�m����+�2�w�Q1�C��]]��^���Eٟ���vR������]�&+�$nID��!�9[?@��	n�]4^�sD��6Ww�G,�grPJ�F�+�������٧������'X�H���RG-o&�]�����i��zxZ�w�[Lb��14Lo�׃^�=#?9|�c�Hr�xC�	��
~e�\d���ˡ�/�F�w����C�'c׏^>�9��&�Y�{�5��%VҾ&8S!g�Y@/��g�g����G�Z6s�]��#$��[��=sU��P��{(�U�}�	>GضΓ�/�)Z��LX��v�m%�S��;�?���<��q���af��ޱ}���T��3��漦U,���Bi9���c�qC��۠]�_�����ᮟ�1�(�T�Ѫ��o"DdT��m'�b�ߪ�KPS�f\�&S�]}rǉ'1�w�8�b�x𜮠�~����'�Q��^<s�U��.��֛�)8�&�ݺ��`��/o-���s� ͛�������b��-��ʨ�0�-�ʟ�z]n�����A�X�Q����wζ���;�z�R�&S)�u��è�+ӝ��#�ozJ-k<��eگ�&�s������u��qs�� 4Iݝ��g���c���"|,8�~Ep@«���;�jpI�W|"����"�~��[�Vs�[�}Y�'��sG��\rN]�(2s����#�I\qL�R�����̹o���:8���d����ͭiP�zϘ����~�q���{Uv*�����L����vB�/�C��$pwI���F�R�;95�sj��1�O��~J���]���V�R:ŘJ��ܮ��yД�f��t��� ��'��&�wE�$lӭ�hc!�&_��C��uW�J�~���%��+�Q�1�6 ���'L�r_��s� �	u�}�ϗ�+bT�@�N�.|�y����}p��>�h��V7����I��k��s����9$�Sp����_{�a5�?u=�/)���Lv��Gy��J�Gv߂T�lk|�P��/����\D�9�~���*�6rC�9D��#݌��O �C̼F���j���āQ3lH�ԚY��b}�����Z������pb��\�3.K����a�c����'� �4_d�g�j�A��+���r-�s�α	�.K�4$t�p��y��e��e�I��C�G���͋�@YB9J�x�6�F.W.��t�.�}\��	iC�8c[@� 1K?���F�� ;(R_�+`ӳ5�� �1%��_�b��Y�m�(�u}|еK�Y���~�g�X⥋r��84��찋��(�[�+�ѷZo޷>D���PG��@(���PqA��ՆM�i�X��J�E8c.Pغ���1U�xñmVm�q�J���V��D,2avޓV�q.��2�f��nZ���KԦθM%�.��H�wuq�C����1_}��8�?R\IȨC�+	�珂WK֑��X��$���9���T�O��l~��|g˾�M�w��^���JŬ��*�ǅd7��>����g�kA,�W)��sв���ύ% ���5N�sV��2�2��,7���QV�LM&b.���Kw>��g$ARg�!P��H:�]oj�?̦չ������\���Կy}kΦ���9��Q�g�8�+$*�����Z���9�*����B%*��-�B��DA?��-AL��g�r6ܩ�2o���)�L�V��g���qu#�]��I��M���u���^!u�	qV�QV��J�Qi�QgۺO G����(�&.��

`�50��0�Du9�2cYgsA/�|�)�;1
a�7�cGK��ahr���v��ŌaU��jaN�x���Y�.��ϟ�}�m��Ο���^�.�CEK��s��DkU ��=�9�`k:M�j&#;g�{9̈́yx��j�ж0��uyR���gv��ߕ&��.��]�B31T�6�@'W2�ӹ��k�
(|o��ʙay�-�j
~������8��3��8x��[��Y���[6�X�yv#�d#gk�L�ws���D�:�\1�-���G����t����a�8�L��Z��� �l�y��A�ʙ��W�q��Tv1 ; $A�w��5~!�%�^S7s즄u����=�J�D��"��;��;nvut�,].$�EM�QΝQ�\%�G�(��6怜�њ�+֣d�ҥ4^h5]+#�H��_UX���o��ew��=Fȡ��T�q�ٙ�A33'�.�.q�p0���?�P�r?lJ�ݡ]��R��?����t(}�H��aOݾ��(4AMd�l�����PA���7��qċ�x>����ء䇂�Xe�M`�l���SI#2H� U�}����ϙ�j�Pr��Z�T��Z<�* �]@g�1����,�/�?96��7x-hRdV$�es����k��4f����={���T	��8�|3sڜ�N
w���_�DV%�A��Y�s�f���}��1X���W�7��DҀ93�iûF��ʄΖ�x�nF��ÊI�vO�l�W�ܝQ@�p6ގpZ�mɖĄA��c��mN���$�B���n <�/� �{��R�k�h��z�n����"{A���#�J�"O{7�:�j��NY��~4�����a��A�y��IoDOV�h��\m�1����ѳ_�5+��@"�t��Zm��[G��o�p$���La@��PRq�Ž�j_�X(�F��BQ,�|���l�y�Z���+���L$�_O]�p�^.$���8��G�si@lUKa.�M�6�����:�����T�sIt; �A�äJ:"J;𹀸�y�#�v�K�Ϣ����h��[�ت��*�� -�WW�(�S�,S��?�e����&�	Q��2%���Qgy?�P}VU�97��RU�Bת�:Y��h'|����HU��R�x�\�/�3���T�7���W>�nig�ǆRl��J�����?_�Bi���ȸ��"�Y$S�4o��	W�"������g?��F�/m��~k,/s��&H�@.�ͨ�����t,-��
��ƴ�JU�T.����[�2���ds:��( g!y�������w���f�1�pb���If�M�}U�B|ݫ�A��Ī�H�qJ���8�5���Z-o��%��$R���U)��޳V|�n����NZ"����`�f���[{H! �S0Xޘ�Ҿ=�?eb�R����;���&�n�G:���y/5X��Ƚ�c}J]m:_�,�/�3j5��C������������=l��4-;]1��[�e#�Tu�������e��6�G.��_z����S��`�:H�>�_���
a�����dڤ��V���d��f���昚�8�<[�7�H��HIE8t������yNtI�gP "k���z�Op=�Æ*�,��)�%��֣�ylSP�	����渵�f���y����r��D�=�}��L&�ݼ��1N�m��'���k���l��ax����S���-�
Ճ-w�<`�UJ�iץO��A���>E�s���D�|�AĆ\	+�#� {R�b��K1#x"�p�p��ES��y��r�]/ct%=�{�(�(�{T~#�k��EM�O�fM��)��9jn�MO���0Fn��]��PA੄A=M��<?$�aΩ��}��+�v����S�p<��Ɲ�&L���YI=�AI��X��:���a#�7��,����7�&�[�c�n�x~�囱U�i�©~��ԃq��<�\�J�J1y	~��·�^v�yr�<;X�*.�y9�o���+�ڕ$�� }n�7�&�Xe��@��P�>� Z��L�Z��@��`HXQ�a�R�gK�6��a<U����7 N����b^�
�B��������I���e�ai\\��ɗ��� 歛Rg�b3>海r�5�v��1�7����N���<�S� o{���ZH�"�D�D�Y�*@:]-sQtݬZ�I�C�F��&�egQ���U���iRb�;�����v�O��2�#@Ba�{��蠤�6�ܥ�BZ�����e�r�������6�p|��8�����|��ҵ�����h�po� �_5�GÞ�'Ѭ���v���%8�g�M��ݑ���m��ۺ)M�2{�KT��O��5�7]n��)��$�[��.z�<�-��㤑��D��Ѵ1 o�w�r҂��*0?y�d���]��c�چ�Z���,��e�!H�p�?��&���0�� y멖D�74���*��L��&�~ht��Ġ�Z�kt�fH5��!i��Ѡ��;�`��; ��Hѝ��a�乔.���~��
|ҩ�K�>�����̵=�=���x&�,�uݎ��Rq6���
8�d�h�<[�2A5p(�v>��o��H̦L���h�p<��6PUv}��`��13���99��A鉵���2��z�Y6<nW�mv�qx �-�*?��5ZN��{+�_H{����d�X�	0C�{3z�Gg#`�����B~:	�v��y�b/#�������
�t=����2H�m˽{qn,�x��B�A�x5CS�4��g��\P�������=Ȣ���7C�_켺��,/[��egq|h	�w q��E�w�G�-��H.6�A�!nyO杉�Yt���vk	�͖���>92(5N�1%����ʮŊt��o�M`�PT��͂L��J4X��D3-���T	K�Dy}g��y�6F���)�7�6h�~��R���2�z3���4�#���վ�ћa7sɅ�)g���w���̮��)��D/ص�L`?�{�N�@�ƈh��BTx#�����������ABm�y�p���q�&Bk�9[��a��W~9d��e.�<D%��� ���`��P-5��&*������מ�y2zVJ�����Ȗva@?/D�Cdshq�M�wk~d6aӞ`+�]�N�H�3`�!w���U��N����'5f�t끥aЧp0�cB�k+J���	i��;f*�6�<e�W�sŎ'� .��wش��.��1bc8k�%�� ���9�|71�}{QD+|UI*$����"�2�6����LrQQf�|���� ��Z_�^ܤ2'�#�:d�?8�1\��U�AWi뭛�v�Q\�;@mq�1�jD3��Z��{���e�����Ƣ�Lx.н���>��<Xz���';��t�0sQ�ᶩ6�s4��4ݎ�Gi��t���J�~�"D�BM��{��2ל,����_��ՑP/4�
�-�	�f�Q��m:5� Yq$�+R)v��%��%;^�+p��*�C���7 �A؀܃�*3���J��JR�2�OG��5A]{����7��y�se!oC5���
�p�N��)�k��A�y�}X�ʐ(�&�nPڰ��T�ǫ�"���i�}w�{w��^�+� Q�P'���2��[r3�$(��:��薖U��ɕ���o슄}�J��9��o�����|y�j��������/Uo�t��{MW����_�����WN�f�����_Cuu�B�mxi#L�9�p?Iξ��Y�Y��e�\��o/L36����&����U���hJ�E,�F?��s��IE3� B-F�f�g��Vy�0&Aml�1ʇk����hv��F� l�;����OtYV�Г���٢�h�Ja�強���R���}�Ն�7��k;%��d�)X�<�ӆ�T����b�h��~׆��;�PE�I3����H�T)MHR�7�z�;ku-���Y�r���>+pU�*�nqV����Y�2bv}���+�U�5�3�1Op��Ng�5����v�q���5kR��E�K�!�OH}7=�Q���U5L�kضp��q�b#�h8�Ra%L"_U�"�?d�)���Fv��ʃ�:������NK<E���0�iR����Z��j83�Zj���Fd`ݯ!���CVv������O]�D�#!��^ ��!��y}
Z;�~7���t�z=�aR�� �*��[�~!������twd�$wa.c���N<t�J�Gh �e�7�,��C�l�����n������[�VP��/��C�R0�4�R�ݪP����E{N�^�I��f�5;���~�'©k�)@Pb���.��\����9��{����]3V�x��?e��w�)���+xi��MYz����b��[�e��-���[v�<����}1&|з,���YUy�%�˶~���t5H�wl_f������!{��]�0)َ�A��ǒ<.J~�PM��	 R/2	`2]Y��������E,w�� �NP��t����Wc�Os!KE!������>Hţ� �.��߹7���H�<� �3=�l������7{@Õ�-����ocTl{[P�~ӔRjQ� �g��Вf��q�}�\3!3u�,eA�F�� 6�j4��cwNQ1�6S��*t��B;����<T��c1,]<ů!����4�hf�����=7���>��+�0΁O ��O����x.u���bj+�� ��s&�Z���k\\�3"� ����z�f�E������Qa�}[��������O��z�����rr����:��lMհ��e|bB��,b�ڜ�N��e
3�6vU}q���y�5t(�X�GX�%�콑��9ӡZ��U��ܛ���P���L������h��.�.e]B�\s�W��7��C��k�#2?�ٌ|�3��x�����%{&Œ�U�1���W�^�{��k���0Cmk*�ٳ�z�p�%4�;��uY�О q�>Ƿ�w��w�Zkވ��x�t�B���MeD����{oG���ψ;q�*6帉w��+&�5�瘖��I���ԊC���������߁.���	�/�h�o��l��۟�NbðJ�����l8��k�J�nǫ�+��޻Ţ�����*X"s8W�nn�	
w��h���9�����b�cF�a6����V�m�!z�6�n�5TG�x�l�wX�,������4ACS5KJP/C��Δ��܏H{��Ԩ5�[�z��q��QS�S�>�*/����[�h���.���}	�В��E]�%\���I�y��z��[�-v��Q�j'��Ǉ@�#��v[&���K�N�{��ދpqh��`��ܸ)<�	��[�ܔ9���ۭz�;?KAi�y|�O�_���gg�lG����xhN��_���B*g]�G�ʓ�a�u}G-���a.��Ұp�d��|CB.�j�U�UP���1�um�y�W��l3��,��s��J\��R���pG���#�xȁh��3�Z��Qdy�O�2b�:�j�j㐾>�q�t~�I����$��f~�I[Q����N�;��ǚu�3�����B ��y��� �?-�K�H���3�hXߺ���0o�.4`�e#��	w���SY��T;������qK��+��/������|����{���]D�Ed�w��(�90�p�i�p�F��r=�3P��-���鉀?�&�Y%��CJ���v�u�%ښ;7����.���1�Y����J�r��k��3��'��P� U�X�	*�ӥ�|.��,�d(�J�X<��?`�m��j%�H�`��p�>���E�ڿ�׵�u��E�d� U�V֮�D-�O�Y��!8������V.�,�Ub�N�ڽoNk,��9��1͕�I��!&5h��~�+f�SB�h�L6ӧ	�N+�ng \hr�`�@i^!�P㤖��Y:gH󧵦@��Cr�k L�	�x%٬�}i�{%�Io	Y}���=8��ٛnqK=[���0ڰ��ǌ�o���"�*�_��֎�O�-4dVɻ�Ξ���0((K�]���;���#|ɰ�{��5�޻��|9�m�����U4z�Z?4���M� �����*Zl˶�����k�K\	0̤Bl�5O�HH�.���e#��%��ȷڔ��d��P�t��55'�$`?����hۆ����� iD?�dpy��.�}X|��^�$a�����Qf���Ǌ��*���2~]R��OM"+���ޚ����T���gyҥSe�; ���VTCC��x���M�[�o2�-��J��;	Kaî�w�O^/9�9s��V^�C�����IRǨÞ��K"5�X��ʺ�=�s�B�l���wu�������[��t�b��8���u,���B� ꙙ$�2#�m�l&pa"�!�檁��J���G�cS������,��	6}�h�\˛�cw��ѻ�����*�t��(^�RF�m*�Ԫ˷�(�;F1���w}���sp ~�	,�q��V�ߺ!_�5y�E5�Je�H��^�t6eL���l�?T*�l��D�ԣ���ږ�&��bY�R�f��ڰ����B��m�&�,��I���������K�G1��Է6��<�;r����p$r�SJ�jڌF�����k�Y>�ުNu��Z�K�eק�c>\?54�UD<�b�I���	�Vx}6^�v�U�������ek(	uB)8����?'ХBf��/��T�G2ܛ�H��H�"����
�ކ/k���Nz߯zW� ߠ&|C5�jZ�e|�h�$$�əٕ����_��Κi�{���Osk�٫x�W�L��)Zw�Ť�I������pQ�*y�̦���~i�5��lN�n��68h��ϯ$��p�b/��T��쇹�ϸW����d��#��SN��B�[2h��C%�ȑW�d�U^�X��W�m�i`������ޗ�9�,'ym�e�KX�e	TdW���~ߊ��o��0������xXF�ݱ\ �2�~|f�z-b%�]X��6-��g"YUd�"G�Օ��u��i6/��e�B�y�<U�xx�b�X���u����E�;�s��3�c�~��/n�Wٿ��u!�E7�<a���^``��H�ٞ�E�^hdvI���C������Q9jW��	��������[��>y���g����}��[�������s�������,BB�I\)	����3�pM��"�Qx��4.'X�
=^��hY�a,���5L����¢^(�o���W��F�j�lj�3��x����/�ǹ�e��e���ӥ���4/F��L*��X�΅�­�������%ו��^_�'�oU*��ACr�IjDp�Uo�����**׀��[���'�j"����w�,�"��D��(4D�E����L��Q�^a�u���k�ڳ�(�ƷZa�c{D	�XsӀ��"�!�%
ZZ���wT'�����86��CEy$��R	]�!di��,ü�qGܯuY�Vʣ`�ѩ�^N<e��ٍ�y1��4ԉ��=����a��`/>D��7vM�B�m�`�tk�R���GKU�+���:7EYl��끾��o���*�EIZ���z1Ȗ�^KcI� ��+��}�Vd�����3pz�C��=�ʐ��z�_B����Z�:�k��lHل.�p8(K��甹��O��_����=���l�`T�a�2�w�b�v�m��0�}0�M�8�'��8N�X��B \�������]��ǆ�۟�d��ED���-[�GJ֙�L��g� �?�D?S�%/U*�Ѷ�:W�Wtm��+�f�UX�/�U�s������k=�(ޢ�ط:j�L&=��&ŏx��e"`� ;�a� ��?�*A�W�=�C�3I=�Ai���n?�&�*=�S,��n���
��4��X����[=K�\k�4]=(o�m�p%�۠��i,���zO&+'�y�~�V`C`VlHT-`��Q�~ۊN�	��z��y�L��4��W#A_Ѩ�ï�9Z��&��ڈ{|��Sf�6����%��X�Z����*�	��M�y��I� �p6�U��g���+��ph�vr�s����W�ݰ�lUVݏ�܂	��8��k�e{��B>3��`e�CQ����}����O<K�3=�ԨO��?�+���j��%���g�s�$�,�C���D����ێU:㛮F7XG�L�����aS]y".v.U�J߫W@-�5�6��'A��͎ZT������wH,�`s�W�ڕT��l����������9
�}(zż~�70,g�w����@!�f�W�[���iSú��p��,x���v7� �YI��.��؇��V�aoEr"�,�U��B����v��^,�]#�3B&�[�@C�2%��c\ia�Q�j��3�����B��%��Ǎl��y�~��|k�M֖�,D�D�6[sPg��7.��~���o�R+�Q�mI;e�4��V�Z�S���1��c��@�s�.>B
.k��)G��Cj�����Y��GFۃb�)M~��J���'i#�/ڋ�}���'���E��	 :�eűM��7�IuG�1�{/����g���P�	m:p�K)=�)�������HqRB��f};L~r�c���*�Pq��X���V�_���i�)��EH�K�Jʱ0�)��:iO��j���{]p�!-)j���ʆB���Ho�~�4�7�kK�')Dy�ȯsK�fږ�ׅ)��Քԃ����9D{?8�6����ʳ	����%��X���=,8:���4�+R&0WB���@�L�(ˆ8"G�������R��J/��nٿ��Tȿi�-r��6Zr���b4��,UL�a�o�	̳TV�A��Rɪ�n�`���#��S���W�7}�q�9ӦO"G������S:�ʦ�^�m�����a��oSJye�Eb�YE�.�6a�1��1��C�tcv��r�kA�Q�ĭ���KT��k��O��J���@d��V,�����n�S�VE��X0c���t�Ϲ����e��@C=�Q��e��j㝗����c��Ƣ`�������#en$�hQ��W+$�q|4���Q��ԃ4ʫ��Bm���ט�ɼkG�r�5g�V�d[	�u�M���@��N���*�o��s�&����F^r"Fb�y��R�X��xS��`��j ��0��0��6�����hB��H�*3�k7k�� �N� �|&�B�Yg:�b|��i� ��\������i�$�3�I�idk���G�,PR�!ۂ�I4?a,�6�(�.hj��~�4ef�������7�Ul�1F�ѵ߻���$���t���h���Hh
�)-�q#���)����`��!�3��ɤ���$�Y��D�����V�Rܔ8xa�J�Ó�����#����"�"B����%�$H>�66'f�Ju��Y/Q��8!ʂ
� _����M#`�jpk��q�b�C���p���Sk>�K��7'�"Vkq��&b� ~�mW\�&PK,f��V�F��
e�ouYt%�Xp?��Y6�TY�N݁b��Y���
X?]яv��ͱ�큛.o��{ 	�N+3ki9Cg��HH���.��V�]��'/7o��FB����{�8 1>�������Xc�(Q�H�e���p�rpuu%l~`ϴ��߰o 1�8�$���q#��]�+U�1~�K�ͧ��tET����QxD�3�:w6@�F��n�I�$C��7��{7KZ��d^����A�9��X�V��h����������R�sxl�0�DF���CPm�
���x��ܚ��KJ�,�|�󋺗z4��&>���� ��VĐ�������̇G����ߜ�9�&��y���P���_
��3�"�K�I!%�LA6s��͑��C�� 戠�KI :�H�ྣ^��+',,�xG��W�������,�(���?H���'o�)����X)�(�1���ܞ�nX-�E�-$T��.K/
��K����uG�S��Wu(&��k̒���E���q�Zq�N�и���ev��ʞ��&�ipy��GG"_�
8���#Y�x�5��7"��
�� ��kx�wv5B,��!M���f ̜���Nm C�f�����[aT`l	",o=������e��N�a���!Xo@����<G�껍.338�߀�����߂�����\�����b�p+Ͳ[w� ���R��|K3 ����h3��N��i�8;�g��q|�ڡ�mKE09��&��l��8_Y4B�n�&�6��m4-�U�>U�B-��CQ�w"5k�Vը�6�FD'��^���|s�.�5_<v1xKC��m����x\�3�w����SW#�U}�c�t��8�������O���`�B�)�^m�y�t�@GA�\��f}�d1�N���I�|Q2��W�3 ���o[���%E) �yܖZ�����OH��{�?::���R%U�|�Y�c�[�ׇ�>|<�t|15e<Q����W	\�/?��=����W��!2,ml���b���!�Eqԍa���6��tK���q+r�80�4�)s~#1��+5�ca5bS�@x�@�L�Y�V�pᚍ9}|M0,��s�S��ަ9P��gG ���5�J���3��'h�����_.ص�m1M���٧S}Za�?E���@4=�́������:;35��wDWM��T�IQ�d6X��[��1�.�c��(`����|`c;9,���o�5�l��ȌP�$�-�0Z���A�Ԇ��Z��������]�2����ߥ����W Ư�hU��ގoh%��D_��{s�t������fSE��u#%
�R�x&����cL�݋��Gn�$�9��r\6��+y�-��c O)�+"=��R8N��[H�\�p���E�߼[�� ��IlY��65�0ވ�Qk���z7M���*γ�9�|�e�B��[)��Ž���R��&�����\/����`8�L�c�6�hCL�1��d�3���I���b49!B�Y�{�ߊ���ϔRɱu���a{��³q�B�|n������M�z����!Λ����ܚ�������%�Z��୞�A�*�(#Z�-�8�'MM�����;�.����C� ��(���	�ն�t9Ӳ�N���u�_����F<���6?��040�m����=DX��D��i�Ֆ1^I�G���ٻ�f%�8g���YY�&2e��/��t�-Rw&��bm$�W]�ϥDЩ���뤃��<5�͊��.n�`�Lץ~��ږ���	�$�sR�|5
]��7:���q��_�������}�@�0�z̦]�����r�d����ÿ��۔��&eƀ��3�i����̹�.�N&�l�Խq��s�-<�.}s͛�5A�w����%�'$���E{ލ���(�(��^F�>|��2Gf��u	�	�z{�gW�	,�M���V��l�
�<�D���S�!J1c�D�8U�Eғ(%�l��.8W��խqɻ�W��q6 �g��H�9�(�TGt���b�;������$�8�!���N<��L�2ͮ�EުŴA>�#����
��.J����"�X�ԗ���V^��=�F�$;`6LP�\z�iQ�j<�[W�����Y\"T1��i'���\�
�sNG �ߺq0Q`����\e�O"�uP=f_F���sR����?7.������c��Z�Jn�"���N�S`	�gQ!9+���+45������ �屙i_|���8���`!p����`b0ج���Q�!&�qJJz�����TͿ/�Or�����	A�d���J�l��-Q�&ۗg��4�?��D&�l�*�#��b�r�dTe��iGϋ�sZ�Mz1��|��5�6<�A �1TJ�#�A%���^'��v�@���.Q�p_?[n�����*[FS�� ��B���
�ö�&^�±�<���������k�oԋ@���I�N`��BP�0�;��/7�M���M�(d������Y���Ⱥ�:j� �hP]�V�)�߷ĩ=�'��vf��l�R'S3�h��t�����Q8�^wOљ.m3SET�f�N,�%��e�!nW�~���΀��:U�Y�Y���)�d
�V�����F�ӥ>/e�6��0Y��s�qT�����
��a��B\q�l%CAǗ7��}��ħ�K�xÄ88l[����C��ƮB�ˊ�dX4�k&43���M��!Zo�f8ˁw��EaymLY9	�.)�M��֦�|uϘ^��/�;�����#6MD��� �Q��7}�P��Y ������!�վ�mtz���4�����L)�=&U���,q��0H�x!Ő�#Y����ޯo�б6Z�N_OxM#T�lG��0��~�T�H5�x�}B##�8���ʙ�Vљ/��3�7l�1�C�t)��7��C�5q/|�YF�h����(����E���1��t����_^fKz�ō�~{T�`��*���)`�p	Q�2Ȳ�l��0H����	2�(�8�a�i۰R�p�[m��l�v�i�mP34Z~Erv���Rf=(c~��Aێ6Cr�9u���VfM�-;��MQB ��:�I�v�/�e�T�@�U�d��8A\'g���2NH���%s��A�Ls"7L�^�B=��RA%@���+
�;@����� <�̈́p�Cam�K"Md��b#&/g0�Sӳx������{i~�}�>�JUs��'�
}�-K�ٙ���[�|���6� y��/Y�˝�7>a��A<Z�S��P�*p�rv����J��^_#98g����0E������o_#��!h�����^�7���Zv�=&$}������c�&M���l+����Ǥ�����>q�@81�f��toĭ8�gw�0~�$;��.���t��7&�8�7����$WI'�X�i�-u�w2xS�f���9%uXJ$%]mT��"C2�ߑZH��^��=����%�ѹ��&�4�)7�u����Kt��~`�o?�0>|�Yɛ&���Ms�u�at�s��+ Xx�Õ��:
��
UFs�J�P+M�8��/�v�{�R��'SYeԳ�6��(�2^Z[��SQ�@��s�o���g�A祿ڈπ�q��Ŧ5!������l�>���o�@�=8���n���f�T�=�
���zϪ[xMr	�){��\��qi�Q=�F��(O��	��T���iW^;e��b���%���`�W���$�s�Ys�U��Nw��ݥ���B-�[��Ț��OF�� P��t4_XW57_J���kuѬ�O��ǰ��1��u���$�[8�^�"�f���1x�o�'})�á���e�0�: D�&�/k�U�j�)c���C�WK�����<�[���luE��d)�"d���/�\g��̦r�׎2�܈慎�0S��𢦲ɡ
�c��Ma�e+)l�%߄�������K���� �2K�=�0}/�r�m����{��	�8�GD���+�R/�B����)�by���T�>�n��`�t��(Gg=bjr�tsצ3wp4��\�^�{h9�{�Yt7|Q�J�U��U�W��� �E��T����q��<2�:�����
����|���?�z8E��/�f,�E���*�θYn�������ڳ�ޙ}�Wg�y�Ӑ[U�O�����,�A��UP��6�@G��lӅ�˵_g�:����U �w��]���Ɵ��@��1��X�u�(C,W���.tz�S-\f��]�O>`g�հ~h�j��<�]����xk�8��UoUȣ�5��U���)=�Pa=�+ ���pl�F#Fc�=ߤ	y�H�\Wo�	�Ҋ�e���e��1��i�Z���L�(j3�I|h-��z�Q'(h���\瞇{���4�߉�~�gX��=hӐ���g�I~@���	D��~G�*C��,o�����GX���,�nyq8�<n�2c=c�S8f���������0����Ik��8��|���)�3�ކ�D�V&��l�t�/�,��U�,*����0y*0Y넎\�����*N
ҍ�z�a�I����׮��1v<��.��/Č��7�L�Ch����1�s�D�Y��?��5�����f���cէFʮ�d>������=�(X�r}��,m��7�#N8ӱ��GB���`�몏zC�3[�n��bB~`�� r��p8�װ6%J�d��*���+=\�|���5�+�4�cy&�f/���dH��N�-���wM�25��e�����y���;�[�G�M8�.Tҧ��r�M<���0x�x����2GbDG�'�%�lS=*���Q?��`�7HM��%Tfݰ�R�"�吏 ��>M�Vd��gR��3��G\���1ͣ՛,�Ȋ!T�K����9���h�`�_쾶t`�fH��N������<�w�r�v�Z���߸E����-3|@���Rh�=I,C	�D[��}d���G�`T���^��� e�Hicwɍ�a�W�)&���NL���Tv��>ma�e�;�x��	��q������ʨZ��ƶ;8�Xw��6R����6 uB���ߊ�&�n�l�v��j��D?���2�i�P�B0#>�nJ��w�#%����;J��V�j��s����%5&JNi��T������݆ UB�3�sf���P�c[gM�S�WF:2Q8u6��Q��|䲦�^���"a���k��`"�P݋=�$�`W�w�]�E��t��>�9����ST�e�ؖ�K��}��/�!$v��W��`fFs�i�TS�A��b�/��uw���Zp ��������jT?SO�-�T@N}@'^���[S">���5w��e��!\Ũ!&G�"�
�	��O�W�g�(�N�V�ΏپTy�,���b��D�~7�6��Ѕcxذ��_G&93��k޶�IjQ	�=G��܃����N���1"�:�z�IK�<��f�:o_��td,#"�R���®T�SuX!^���[6����0��*����HS:��jQ��k��$��E��M"8�բ�T�I�[��IOJ���v���JJ��F}\���ƁR뽕~�W�����<7ݐ  �h�NbӪ�_ ��f�N+$KHA���
���-���;D�n� 8/���>#oJd�a^G���I;		��%b��~+�g���: �oMN�,���]��B&�Ų���cч[ 4���335thY�`�B��4O�g�p�Z_�s_<lM2oǲ{yH�r,�i?���c�f��wrF��v���I+t��慛K�-��xy��(K�Ɲat3w�+�v� �d^͹p��*3�f%T�L�T!��5n,�s��T!��&ʵ�!{�:����e���ߥ�:5����I�kmh)#�k�i�a�cY�zĎ�ꉛ���bة��ڝ�W�y�
^�sɷBI���B<{$�y��uT��
�C�)�-���W�h�d+2�l�r����ğn������5��Nb���Ծ�$���YD�X$P���ѫ7�+F3����KG�?c,��=���� �D������S���8��h;�V��'ݱ�6��s�b�_!� Y$H ���^=�ZI�U.�k���pCj���}�
��}�qm�k���Ӏ�ؚxk��H�%GȨ��t(�|��d�Y�*��ˢ��c��N�)��"�l.9��MR���t�};<2�_㑊�4ȻK��[/{�Y@��Q!�%2b=�d(Q�� ��{��,+v�a�k��'���#��:+��ʊ��.��g��c>�_���4d4���l�ʤM,1rX$�щ��S�Ǔ�fLOn!��!?�]�T�L_p�,�B�va�)�$��@I8�G���Y(�dӴD>|&\3ƏJg~��r��Q�ͻ� 9i�!��<:ʩJ����e۰\];���FJ��~�6�L�tڇ�� ���@�8X$Z�:P�MT2&��hf��j���ܐ�8s�y�ʔI�b�;7�l����4���z��ۅ��tt߆&G�a�-2�@s	Ѥb���bPI�+*�㵪�����|Gϴ�)�@oN|c��(�B-���״�����#U�7���1�{�@���;{�v�?-�:�P+!w�[��i�ɫP��
a�$�w��8����514M�4,�V���XX&}�Ï�sJŕ�6�$X2��d����]B��l�d_?;���x�>\�ڭ[�$Mc�:�%��}\�@����TY��	Y����h~>����8_U�&�Xzӿ*���4$7,���b�Z����.Qp�Z�\�>'!��,UP��|����B��S�Q*�P���m�P�t��'��xGbIa��)�5=g}���r��Ra���;5��*�I�`j��X�k���p���gU6�"q�Z�_ZbN״ЀR�Ǝ�1I�=BxB)�N�ꔉj�`���PRQ�����Ҽ��3���9C`0^;��~>{�&�m�\o��r��Ӣ���5uT`�I[+��<M�6��L-�F<g��m^y�
UuԮux=J��7]��Ct�d�W	��!�{���f/�	䷢�;��-�>�m)ħ�h�O���PnV���g_� �� T�T�|7ZZ�ń�2�LN+�!�W���d�Q|J����f�g6���AV��-NABE��Ѣ8���L�	�M�t���z��욆�;�*��yS+@b��o�1Y��j��	#GUjd�����O�R�D�K�+v�Ν��е���?/%&I��;b���^��m��`٬��n�՛|�M����5�-�+"Wt c'd �-�\Iu���J�:�7�D;ܪa+�	�{a���)�j9�d��z<l��AD����@秊�=l�W:�p
���Μz`]������]�K������t��~^;A&{pO�m���},|�S�� w�|m�����@��w���ɐI*Ax3Rޕw��@���;�*��kx.8[�RZ���k(��q�2����r�M<�����8�<8;~=��l�r���m��p!��%P�a��i�c�ҙ#vofG����7��3m��@a�(��B
�U����F�$��,>�֐[ZU}���Yj�.���M�3����� n�s�(!C���ۆ2v����W���53���,؏SE��X��|��G\U���$����� ����6��>�D paO�͐�bh/���`��d���S=^BYJ������8��dġw3I�i~�`	Ja���<j|����1��wy�+�܉z�J9l���3����\��?�A՛d�ڎ��J��O�E�A����J����_r����º/]䬄˃�Cgb���=� �A�X��z�_$g��+	�,s6��L�%%�y\`�6�ta}� \+�������&	+ٸ�gT��H�Y\~}W1�F�u�N��<?�7��֯������e�8I�<�)��ۜ��_���k��@� ��J��H�ݛ�c��ۤ�#) ���'�b�CZ�\��h%������]��IDmnۣ+(�DmX:�ΚM�AT�u�Uvcكh#�&
�C[o��H�|�#[��e�:��S��4'x7W~'��{��~��ڔ5j���qfT�����r���~��z��}\�'��k<��|
�"�-rukUqnd���)lg��N
���4#';%	��2>���	<�Nz�Oej��^���-g�\����\�
s���4���;�p���d�ꋺ�T\"�t���"�j ��-b=D#�Jt��[�G]B���˲ϕ_Ae�#OV7�kU��}����$�{��<���-���-z U��h@���*u��_�L0*�C��2�6_�&G�Ty�����(���?t��^X����W"k䦠g���b�
ͫ��b񩌚��( ݢ�*C���S"�}^��n^��TD�s]+k{��4)���E����D �qlݘ�p]��
�4��R�C�*
J��S�+tL��}��=A�l��v=�ko�_���G����-�bI��!�z3(���0v�l��(��v�AY~�sFi���ż�,�,̹$�)}3:Xnd��3�1�&�A��g�M*��W�Xܼ�l}�R�n����P[&�+ q���u�[�&����b���۴��m�}4<�4Ĵp�|���*L�j���pJ���~c�5�8�NCV�!���h�h��A���x������+����T����t�J1A][���T� �w��o�_��}�"B�-f���\'ؚ������W�69c2��9���m���'�i�A?̵��k�J�y!���P*Nf4B)	����b$�xrw�dz"�y�C3%٦�&u����@z�N����n�{xql~+�T eX�������f�8X�� �J�%��P�x�(e��Q+�J0�(-�p��ט�`0LG��l�8$���f���,5U�{Ǌ�I%rx`a����	
�~j{D���@��_hZ��r�`�Z
�y��38-��U����=�U�t�Dg�}��$H��3���Ïsm棟ԁ_����E��wZ̡kfD�b�W�'9��1���CQ����I��aV��y���u0�=����9���'����Py��L�%	�a?~.Td�e`�;�M�Mr���ӥ��HIX11Z`N�;������������d��!�6�M�����fof���Pڀ&��%�fI����1%a�fT�Щo򭯡ɟP��0D�j$�T���(l��V6� ��Х��j���c��
�)ݡ�O�f��)�)ۡ�~4zCT��ct��w/Х��IF����Ƽ�!�gΔb#&&���$
�WCF�®����uɁ��I�u���^�r��y��o�U�һBܮ�,�a��J������]u�V�K<x�H���Ħc�|���y����3X�iv�s�C�6���Gr���n�]����[`��GYF��B� H;.ہ
�ED�-'a�:l^���+��&�M��"���`|̈́I�|��6
Od�L��T��F_IL�����3����W���Y�XẁN"�	�T�&�<��k8��-Gٗ���'"���YovkH�>�W���\�@x�b�^����:�qT)�Ֆ}���he�+!�A#��_�/��2� Q<���dI��}.Ӑխm�l�x���l��b�urc���U�lU��q���{��� }҈a8w�Qn����`��_�U����A��j,O!�#Œ���xp�?c�LH�����d�jP��!4�nI0fӀ�_�Βp�S�?����jj�PX��L\��
G�v^�]VrF�����Я@S�\e��̻��GA0ݼ��L�l4w�V�i�>[ ���8)jL	;��z�o �]�]bAi�ҿ���ݷ�:,�BՉ���x��U;����-��d�ͯ��R/�V�H�M��t	s�+�G�C��aZ	��zeP�_E`����ؗ��mXې8�L��`���{�a�n�ږ�$��U�Kf����<���٢�
�?r(�k��ǜ�^�p��ET�Lm�*�k\}���vz�_~�g�z[[������^�����P���@�64���C���34�ȭ�5d�5H�C���	I��x��\I�RiS��ʳ{���b��!V��Q����
�_��h�-���SU�(��1�G���d���Wrr`��A��u����+�2C��j;9�!'�!F$#�z�p�X����Q����� �f�P
�#}�h�?�_̭ʫ�y?ԇ:�TלPᾪ�}��l̈L>��/A_��NԶ�"H�.���4��ְ����T��`x���z�Oj7���o�J!%�YK��?t	�ųfQ+<u�[UQ�r����8$��=&� ��<aZ�F��y��|;�E^��q�L�fX]DK�9u���D� ��c*�<���Q����R_�"�д�?L��=+��ik$9���<�#bj�\]�WI��!dv��Í�9u��'�h�傢�����5�����r�b0�K�ˤ���3����+� �xqb��U�/�h���[��U0M/�\5�I�$y]Z��I;$0I����:�3��y��G��J����s�*	�\O�؀�U<�l�&�������#os�JL��;�%񏽲��`�T����o���sAh 1�j���	��ơĬ\���x�d��B*x-a�����C����@1�&���sx�̌ikn	"�v������|D;M,#w���2���ͣ��n���Jao�j��ps��7S�\��h5��.�����F����Iw�-��v,�P��h���W/����{��3r9쏋$)�v	 u�R�4hZr�GV`X�&f�R>�5 xd�>ǎ��.b!q���bx�7��Ԕ��5-��
_gҫ�WE,Y��C �x�V�c��V�.�岢�8)䋬�����4՟��؉G��7���5M��ު=�����vа��TbP�b�q˜.��v�%hE���d����_j���4��>����,1�����ee~��	��&�l���G]�3'[�b�z�������c��!	c���7��hm�1�?����%yˀ)��Pq>cS���M�/��<��v���ok$�6�	������ғ�;sf9�-U�AvV�_���&κ�9��Tol3\����C�BA'{/�>}z~7>ν'4�y]�A��ϧ,�Nʵ*]����������H��xk�%yE>�勷 "v������x)]۰�� �?�;bac&*�@ın���K<ɏ�������6Kk9��H-���eK�1||V���ب��FCv��Lڟd&Dc�j1S1���v1k��<TEF��{z���8t <�аq��@Zv���]d���b	5�� Ϩ���%�A�V��E1ܟc�� P�=��&øQ�ێu��+1QS$�e{�&T�eӪ�@E��;���ҍ�fv�*�����	.$z|5����{�B�*�/>�-�b�E��.����	��$=D��F>�w�<�g �{������xP���.�xz��#�Ꞙ�2X��~���N��G��|�تLq���ߧS���h=����^!;��MI�E~�����ˏ�ą��IXK��jS��q�m�X$�~�E䠸3�~��̗p��ifh��,��s�*T�P�=��T�N��z&�ݯ��J�j����uqLDiG�:Դ��ԛ�5Z�Y��k:��}�~zz-X�~j��,q�='
�����6��E"�=�%���8C;LvW�(��A� ����&^M�F<H�$o�Ǉ��-A��T< �<��,%�I��u)+�f� �Α�3�nR�Nȳ�shڟI�H8) K�"~�h�b�RJIKU�(�x�vR"�H�z6P^\�[��k�:��6������LΗ��۞�Ý�*| �A��u����
�8�yV���khr�0��c%��*������U8�h�+����U03g,�Dra����~�w�k�����:��|�J�5��P_���ശ�Dqgb���t�N7����R0�]�����f�L�.9y�M��qI2��7n��h,fH>�;���T���2 ��fݤ�V�D/�*���C��T�%���{�V෉��c�`�%Ol;�_	N�đ���^�,�eɗ�oOH�@�u���E4I'�(���/Y�͕3{98��cd�+ĎbUт�1��{S(����d3�a�js=g���HQa��g�߽��m���~�x�І��E��C��l_�V?����TW���Ͼ�;��M9$.Mq3��zܣI����jYMK��,�յ)7�f���
.��Ѥ�P읚�ғJd�}7@�Ln�TT�.IV>>M@hWk�=�}G�%�$7�� mDM�x"&:Ge	����Ԙz��� 7O�[LB�p��n%�%�⃉	�s�6����߈a᎞u�f`^ͪn��-�v-S�wT;�H-�]�jJ�����ŤR3�K�=�x]�z�����Ma{B=RΒM9�ǵ-��9�ʈ�:A�eQ?}���1��4[?s�Ua7,k�RO�ޯ�:m�c�%����HY�:�2��s�;����g#ƭ7
��������V�;Da"p�7/��`���~=�1�(1�+�q�5Z�����U��D�*�_U
�=�1W�!���\�	�#��CW�
�C�#���5� �kijT$�6XA
�$W���z�<�ng%��wȍ�۝�x��/���~�)�޲�:�� #3�Y^�ogl�n&sn
��A}�1�V�;F�:���5�����V!���p���g�(q�߂B�B�ݪ��,Y����x���Us(�@��k�l�o��r������'��_�:�c�k}�r�'Q&��q��'��q*z.�^|��O#�X߮.�	+��~���/d%�������p)j���O��/��Vp�5荭Ӕ��G�n��!]���6f�҂���f�:�rh�"K�O.3��K����6�����`ݞ��g'�J)���a���l p�2�������RI;V��Q�w����ڢ��ʧ�	|�8���Kk�U`�/�>]�������~u�e�1�r�/T2'�)--Пϊ��o��Q�� I=p�}�:[?�����+�&��*A,G��G~935O��o7��m|�*�{�@y?*���BNx��4���Uʫ�N���"ϕ�BG��W��|E�7
�ץ���2<�	�=��y;�R�bѺY�D�{�l�G�D-�-���w+��3߿B�#�������4����(�p�W�(�d�"ؕ���7��u)߀4�"O��#���f/��� �G?�+Km����\�Y&� �n�����l�WB܈�$�&���!,��S�O6�*q;�iQh"��!LJ����){d�]��M�v�b�yO���$��u�������,m$�EO�UtmC��J���9��2�O)T8����Q�hmb`�g���y8���#~��26�ѡ���Cz��t~�ge���ͽ� !�È�5<��L����=�W��W>M��B���w�>o��m@�̵C�����,�	gw�){OH*� ��Z��;���O�x`��lYJ\�����S�$bz���Mlw��� �,ehD�g:m�\��OW|��RR �%SNM�!3�)��\���L���o�M��Y;G理2�0�Q�4!D�M��Ӓ��>�k������0�8Z9<����"��d�-\�'�00����8�K��n��Wt�X�덲�{��j���s�)k��{s|�G 0ҳF��P=-ʳ�~ho䬎"`i�̌P�p.zcST��%����DFS��!c��Y�K�I>f�؄�L�X��d�+�hsK��@"��i�4�(�R�#�h�I��9C<L��n����$�;��l�K�u?s���ah^�F��?��ό���#E�0��Vy����zƧlê^G4��
%���S�C�x�8Y�x�F��{��ʿ������#ɬ*6J��`�N����:I��1��-�c'�$*�	���x����)%ش�No��:AY��0�[r[׺��Q��!�7hU]�d��J��@����ݝ��B(���I�Y�	�`�.U�*�H��]���S9��?V�����$.J�$k��Pe]�h��T9yi
L�55H� �,�p�&���PyM=�6�p���׻��o�p�i-���T_�7��<�8�h0��i�n_?��������{v����Y�^�Q= N�w	�qk���c���f�1������-���k���;Y�!���V2)��IS��Hے&��	����{���|��R
�u��mS�l#)c���B;p��Q[r@��F5�e%_l�!�����FE�d��	��Oz��>z��5��lR��|�{LT�*\_�^��č]��4�t���)��{fۂG����fü�j��< Ûs{��K5�/=W��	z�yWC�P*݂��	����� K��u���M$���RG:Y��a�M4c��ED�a$���VZOxm֌ϓX������Xό>}n�_�io��f�D����M#�
�*+��!r~<s���!�-hE�wz��\2�R�j�g��<`�rP�wt-~���Je�C��o�-�J�`��፠�d6�� ��p�߼�9~�"\s3wF�CN���X(P�ֽHa��,���^���7��đ�̂��+�[[� �</.7�Ǳ���)��2'_҈�g�
��[c�Kvh6g>\�T�xG���סA��=:b�5�&�����m�5����C�ǟֆ�N�cA����c� 9�BXJ.$Oq��`�|0���_�W�]��X���md�2s��R�a2<֥e �J?d^������=�?)O��Y�ɳS��Ԗ��S���{,Z
�R�w�n�,[��aU܊�˿��q6'���L�Ł�f�T���ʕ��p�i�6j�����OT�Q�p�0�� b��NoX����.x24�P)�^O�`4�7-���8��刾��f5�`��v��ۃp�ҤGx�$WF
. W���ܠ�g�*��{�(p�j�w��y0�|f���@j�m?� {�m�	�1Y��(� c��7G*���ͻ�܀Vϲ�/�"�Ϯ �꼳R��U���*M]�P.[�S�^��� Ȋvpz+^������_Û;���R��Lnɬ踐�d2�rwg��Y:kl��� ��D�M1�c�� Pd�m�Sa|�G��:g���Q�B�T�|��c׭�u
l��������a�q$�s�jt�5�u�|X����l��U�>/���n{�!l�̥��N~y�o��?��@^LN
���Vx]�ab2Z��y���w��E&<D�]O0�VaX}S�s����*���o~�Q���u3l�{��s�7��<ϩuZ���w��t��4��7�=4C����?m!v%C�B��x6I^�d��
�ڂ"车Y`;���@�,�?G�2���FX�yu�>r�L�o��Sx6��6w�fy���2=�Y��g��
�$&ʆ�Q(�x��7���\����3=ܧ������#l���ǲ�ԋ�"̡lֿ�V\��H���T�k� �Q�G��Ԃ�.#^˫d�<��E'���s���Ũ���_��E���:��~3��y��N�s����o�3�o��4A8Idi���ϟJ0r�ds+lp�B���i $�B�q��X_ߐ@K_N��U��7X�5n8u�a�u N5����H­��Y��D�۝�Db6U�܄�2���]��\#���D Uvw�
�U����y3����rT�d��+P�s�V��n�&�@x��h~�V���ʽl|lgaH������e*�'�>�i�3�j��!<�1¼HEE�Qɱ���Rs�62�]sm�l�-��dO���@:��t�6���;��>����^���*����OZ�ˍW����}>SIt]�1H,ib4�3ty���#��~՗i�V��5b��]{��dQYq`���H�'�ݪ���4�Ie����m���.؉,�ĹJ��*�YZ�}�ד�7JLĎ- �a�?Kzé%`�+hByE쟀����'���f��X�k7~���%�ǡ�f����)\��s�pp�J��=6u� w�|b�@��G���<���������pqc�Z�x5�Sq��(�����l&Z<�ģ�E�d*$��7��x�3Y~T*h�u����?ˤ��?��O���)���4?GPr�-+o\�O��[�_�� ��S�gi0�
&�'@��z/kr[�)��BZ�娣�Gj���wY,�,��[�G]@?pg��֟��s��n�'��8�5Rp�tK`I�x�S7?�v��7Z�*�X ����Q@��󕯓m�A8���,S㏘��e^�_K�J�6Ά�� ���)N��'_nɌ�1�rI��mp�8x�;!��jG�#��!VSeʣ��6��B���#���]ؒJz��	�%��m�q��bs=��0b���ÄI:��	t\z|Р)G`�ĴF�����TՍ ��ޡ�w�N3���u$x�*�x����q�ayxds�ұ�Տ��N�w��FJ�d�bw�F��L�p0 {;�.�(�\���62��FY�}�St�3"ׅ:��L��G��[	1����D�١�mĢ���OpX'�}��P{�M�j
Q����i�����)�f⦦n;s�/0{�PN�HM� ���������9�rg��VN���b3�Cs�Q_�s6Cvp��'�$��~<J��c�1^e��P��U��AH��#R�0]4�h^��D҃���x�1w]��� �\�ܑ�HF��Ym�OƜ=�Ɉr+����D�#3a��	ǖ*��U�L��?�8�=)x�ETC�Xa7���s",�v�}c}�ƣ�,�z
���.��_M}�9���B����4�xF��2֢*�9vm��nekH�h���v,�#
�	>.7�� n�m���t�<���0%�$�0ݘ�ۨ��{�9��*A���Y9�YUS]�� 9ݟ+���\@��gN��(�~���XP��l�������Yk�)��+;"T��i������]���/�1���DIq��wfՁ���� �]̢R}��^}��@YlU6;�Bh1�O������ZG�5���k����ЅKr����=�&�#�n%۽(��W�!鷓�J��@�Ջ	]BF?�.�fA��@��/�vP�'~��S>����i���V��"r������(���a����3�򂅆�w2��ӧ5����}yH�.��JΠu^c^
�����L�Ė������P������rQ]�P�[��?��*9!e��o�G5*�'�g����{�Y���=N��~�=� �Z�����Z�ԓC�����e�����_�Y�'%��V�r���(D��D�ĺ��z'X
����X��w]��%2�@���$��4;0��1��݆�
�&�k$���U�d2���ҋ��-�IlZ� �E��c�n�����]2�TS%	��CuTw�Rf�u�ǯT��Y���D��\]�j_NF.aD[�}y�Ĭ���1z�8��L�Y��o��*�."!)�$h�O�oL< �q��YKE3VQM���dFn��qW�"���{�[E�2�g�v?zH4�''��# :�F�S�X+���)ҭ0��.\�6�&x��ɔ df..�Ǡ��g����Z˷s�-뀭s+�U&��)�s?�r��
���!���F!�"�Q8�Ϧ'�u����A�`@���E������~B��
��L�U�!�^C�Kyjv-���L]t�8�稅�oA��誛1��V��ﬔ�ˆ4����a��N�H�I�Z�;�,�ݴ�����;(���WqO���r���0��TB��'��&�����o���G�/)�@�f��\X����������>k�ׅ͌�C\�ܱ{o�[�D���Ɨ)v�J�g�֩/�HMK��i��1t��O9�о;�q4!��뢓��8�T�����2�\�F0��*A�8�V �z�:�{�M�_���{U}1�x;zs��I�|.O�٫���C�N�D�ȸ���	ɴ9���N�M$d����;5lwt�~mO넗�Q�+i��6Ѓt{�K����%������c{�_����e'�a�37Z���`_z�'��3���q�+�bp�q6�kP=]E���39��hJӄH3Ę�Gv��X�U������Gi�r�*b�U�ؖ*ZR�T"�ZY����W`��?�̫`�W�/>�e�q����v�<�î�3�	z���s���CA6~�V1]e��9�H�ש��<}�jo&���z�ev�<�Q�DCM�qoYƆh����e�Up���ڧ\��10��Ūю �g1�kL0��D�^_�x�>E��,�)a�b�-��H1 ����S6���H��R������!��O��N�	C�[tjR_P�$�z�	 ����W�s�0��;\UA�M���H��qXzIa������",F��ܻ�=��|H�p�I�)�ܧ}�v�L�D���2�vG���z|��pB���q��&����C�g0���Uo�N���j+d!uS�N��t��h�&�:_��&�Oy����"�F��4%��?�O���b�*ҕ˶#"�9z)nPΓ�������uJxo�G���T�����oD3�9U~����rY�GIa�:�4�(�����O  Vq����~pz��2���Yŀ�|V�f��Bv�`7�����7c)�moyi��chKEzAh�><���[��o�2��a��׸2�P1C�_�G�!Z8m�#�U�z���+�N �`W�(٠�G��8䰨�A��R��v�*��_�$�Q���A�=��n�x��Y�@����Lc��k�\���4ڿ�N��?� k_3�,̺�3U�M&�e�e����&��eCM��ˀO��2�1y����m�������l�?��P�K�d�q�j���|ɍ�7ŧ��:K��+@��;��I]�����f��5l��z}ki���#��0֏.������Q���S��>D����3���EB�B<�U�TJ����)c�ʯ��w�'��ڴ�Ce��-C8^�����g^F����T�� �yW�&��pà�����.��P��O�Z.qp1X6�e���e�����
��FqO1v;J__��0E���ǻ}5��B�+lř'�1^W{76�:v��I=̡�a���s3�8��[44�'��3���em�aA���0W�����D��3����M�U��f2/?�\���IE�,3�cc*��T42jј� ��P�WTn��M�p�ޯ��W�yMhU,��������ˤ�4]DS+�֠^��U��$���>S�2�Lp�H�I��yd�=��&~�ڼ��D�*b�k��`���u83��������rp�G5)�g�xu#�� ���')��Ř��1\bj�\�?�*�&����6T;�,L�=�4�}����~j0�ԗa����wⷜ����at<끗B�ޒ�Yك&��o*nO�^S��:�v�e�C��`ԉ����n�ӿj�y�[� c*�{��A���p]1E���_����r�Ĳ��:=��	������"J/
zts	���R,�0����Jk���*����\�V'z�|�#�s',��B��C���%00'h.�qY�\}";�����֟2l��!I��ς�lK�kG~�"j�i�E1�q�bZ+o����e1/F9�B2�5� (P%}F�n�(��uH�z\s����})���"}���,su��-�@7��"�H@e3ip��I)Qˡb�p��7�+XE���EWyV0^���Z[]� �	�������F��E+��Hv����SnBE���S߉�L��N�!�o�p(s-TE:���'�(�����~�#{lP����)|���ڥ�i�&�gI��֠�	�ٶ�a�U��?��y�BFV�@����;�
fv��)\Z��Mt���C�s����X8�k�[�}�^�$���3]�X�k�3;�+�� V{k����� �N�y3!s=�(�Uh���YԌ,^M�:{���pt}�G �9����܃S���#�٤��i�b�pp����.,������dDf�I�}5�������.�W���ɬ�r���x���B�?�#s�@ :]x�>[Ӎk-4���T)��q�ݫsC���?є�7Ka�n�f��aD1���4/2k�wQv��}����*��	�xt;mE�ǔ.|�~�F&�"x����3$��(��=���q`��Ϣr���:���
h�^��0mpa�s��/���/4>J1<�U�;�T_ �g;�5�~q����j���t��p���$�������I�K"�Q,�R}j�9椝"��!�#�c�	*N�]������t��긍 �~��ү�����l)����u�=o0X����-�٨��-u3_�	���8H�|*Ӑi2�h(~�����Z���H���s��"�C��u�1Wo�[���3��M{EI�9�Wg���SM&��+,�)2輄��0��=���� ��I��e�[-����c b��TC#���Js����)�ܥ��A�N6�$��{�����0�����7`�9�<,a�mW�߯2`v��O�TI'����1Fx�4�[{���xN"_;�<R�a
`.:�	P���&��|�_��H�:�HL~cܡGb����{\�]�"9��	�%�����C�=�I��mC�0ODc�6lB`�#��Bq����KB�1F�z�rM|ƋpG;����p4��9������#�:`�*G���8(Y?n��]��rl2@�*6������y�Y�"�l��UD02X^"��¨5<EO�F��?�ں���9��,�",Rc_��sK݉��t�2ͻ���U#�T4!���kN��%��E�ֳG�;@�_�3�/��
#a_)��jY�P�J-����ք�<�R[\��},�N�Ԙ�Nlə����A[h���k��r�����Aj�c8Lf�)&�'�W|��-�x�	������.�N�er���_$D�wm=��Ec��i���eR�~�u�3�A���rJ��*�tǒ�쨦� ��Y�����:�5,��S�U-}Y����J�G��s�,�&�����2^6���5��l(�?`��Kɛ�(��L��*$�����j�m:M��w�g��{�}ض5,R��]�}\n$3���޷��]�;	m
�Z�,Wj�Ԙ����-r��u��ej�]Êr��t��� I���l�y�� ��| z�k����2f��'O���8* ��A�ń�?�c�v?|�H��6 ��F/v��c�q�im����iOY�T�������~Z���xv�������/�������FfT(���o�	�֓�M/�G��t\����m4�+�lMqy]C�d��8Ŏ�Ø�����(�������Lֈ~�m��sy�v;��I����C<�ޥ?n�U��W@����0Yƅ�a���'c��p�z��O��98��O�糗�;=a`���(�YT���VmQ�,Q}���Ƞ�㸶5���u�ja�9K�)�����v�����w�K����:�ؓ�h����
�l�h:�/��/ޟG=<�	XȆ>���L���G��n
�o�V�}�Nq���
@�U�CV��H�a	�_��n(�y �%ę�%�?X��`	@��'"��Rl,t�>��A��0՟~�"���_���e=.g$���^w��^��������˚ԡ���|v���;�}����2����s��O���ܨ��f��:.�Ø{"����'�LQ�M?6��0[�s5���i2Dx�}y`����흙S
QĘ�R���L����`���B���] Irl�a��aW�ǌ���ٿ���?��>�c�CW�AiR��,.��Ќ�Z�~�.��.9�̢l������?����;-��@���Ě�+TQ�5>BW�v:m�WQ�6�XF=���޶d;��O�g]8�|r%�A��@��P��K�ڿv��?B�ز��K^�䵝�@d�{���8j�0�Q�+���,ˮ����
�H�����H��ǉIZ}�t��'WI���P:�j�u(-�fhC�v=i-O�'ó}��f|E�G�������?���&��n姹2bś��
�2<6���u~>�$�]�iGr�QVӽv��:|!�5
��J(�B0����5
��I�3*JR�������:tmƥ	��x����� �5�I��]��CX�c"�R^N7U�@V��)99��GIZ �U	���\.�/^1ٹG���������d��!��o@D�v�,�d3�ff���NB;X!�ٽ ���0��-����_~�W��c����p��M�.�!����~���&���@����;�_X}G�0�������s��8���"����0þ�'Ջu��AVdWu;�3�y�x�g�3W]�'aEn���=t?��H	f��T���lk{Կ��4���*a#�"t���'�>m4�;k�P�({�=j+<�I�p�ϽX�i�e�a�-���`sUF��=`h�SY��KԇSO���C�i47*�����Y�R�h=�1c˞&�彾��b~���T�k�2����D�%t�5}���ܼ@SU*�I}�r\������2d6��ވ/�¤�'������Z��;>��2{5�\��m��#Y�y�?�Q�E���Q="��  �Gg��Z��7�=��ܗ�1�RT���?g�q9���9��YKc���}�v5�BPv���Q�fX�T1�����Kz��:q�/.3�4^�JYm��Ty���%u9D��")���$;��m?����p���4StY,3\�����	7�������b �6�,� �����Y���4�)�s�MM��T<S8/�:�#q#����[�מ�?M>�p�fh�v�x���$Qn)ּ�=����)�ݓ?F��c����nM���YYjI��7�V\�8����'w�@��5���Dwȹ��� ���T+8(U�a�xW��s�b�$mU���Lyѯ���e?�᝭3��~L[�qH�
yg��4\|��<RI�����C,�`6�*�F�5䧻ЄH^�9���&�^+5������,Q #Pa��[��;!�=_��B�@��g[tx��	��RU9-k�ךM��nu���� qe�-�@M.�_Q4��v�|�Ձ�G�WT���nu@������!������0wFx'�@��ځ��5�4�RT�C�=��b)*�=?��.L��6��3M@פ�`�h�ڷ�[��H�#^�����?��0������׎���'�0��NOOǝ��DM.TE��6���h+���:�sw�/`j��n�|/Pү$��T"����x� z�ԟ���O����ri�C�-���Y�3w�� RgͥHo�WN���Ss��\�p\�S(F�5_Mnx�D[-�-E}s-�TN�'v�CS11i:yoq%Rlc;�G&�(�E���M��F=�җ������$
��qq1ǿ�ETvn�j�f��[���d	钴�p@kj���b"�bCB6��_��r�9�������M�9�VP��!��]���� ���ˀ�����X��^uJ�`V���;�MȒ� rcL��|"|�=~����2�k��O5�J����o�k����;�<���V̻�&��_%K�^�+������N�i[\�܍4w[�v"�C ��Q� �M�X��&U�W�E�L�3R���C_e6C*�$1�.��:d�#��a�c	�H�څ��݀�4�W׹��x�7:QYg�O��el5up/_�XK���(u�\��s�`��H�� -��+-���0�+���H]�dA�sW��g�	�N���n�t1[�!�>l���MgX@�q{=�7%�Y�ʩw���A��
-����j)�߃ Ke�s'4^p����>"">��E�h��}g�闋�� �6j0��4��e���<�}bZ�5
Mf�uʵ}�)Ȃ���C���W��Y��
�W��� Lb����Ȱ��-cA\w���W�rGv$�Fa���+-g���ȏw\Jgl�Oi�.����Gnl'2m�-���E(�h���F�Xn(˫����w/�$ F:nޓ]�!f���ލ��<Cϥ�m�r� A2�8;���^�%���z�]�;�%zOZbǐ|���Ht��ujHi�,����T�פ���R�@�.��xe�.���xᴞ��~�����j��"����\�=x��[D[��؉�wr�.ӌ���U��K��%9�CE� �V���M	X?�L�P���/�='Uŗv�L�\�{qE���*�IRS��-�ƽ�F�"x�`����S�l4� �^���x�x���	�A3�r�ow�LIܾꢟ��(�W&�;d�^q��`�)�꺆�/$��A�9�t���G,�jf5��Ly�������/��mA9�}�iTԄ�vT�G]��I���Z��L��?�F�p�	0Rd��e�祐�;Dm�E��P
��|�F�4�~[�sX�N`�.r��6Ux�uˡ�p�%�?�FL�D���X�����3fm $�x�2%�=��_�.�#SQ;��T���7�Qz���S�� �Hy���2qL�.%��~5��R�����n9��ڝ]��yR5���gwm���|?�)$a�+��9oʯ_�)� ��~�ݔ��]`�Y�x������A9Ӛ��qU�8�,���f��u�TӦ�����u@fs���+��$Z�����m)2/g���)"$�ʈ��u����_�݁���YV��`ֿ�UlP�����Z��3a:��\���|�l:J&��|�fxH>�¨��ڀ�:���*�f�i��x�U&p���T����Vy��Y�����D��'��m�"��q}`<�E0e"(,⑁L7��8A�ӂ 1ۋK#�:L�5n���w��0>�D����]��n@@����m��?M��:��n4�փ?�4'�V�A�����������A�u	w!��ݵQ�?%�6=�+����U���icG,�g�t�������"��]�*�V �R]!�[�����w��˚'TkY�n~�R��%�x$Q l���c��q��Lpl1֘���0yeq�����tH����梕�AF�Z���m��(�%W�����y\�,pӕfb�=���0�"��ag��,��J)�/:��m�j@�V�0q��p����k?�P'*Io��Ջ�<'1�᥊%F�v=�r���,�-��^?/:A������:�bi���by����vk��[0�iG��Ӡ��p�V*�@�n����(�z7�~;�Td����|s`?@b9�̄��տ�MaHE��E�=�Fz����Sc�aꨫ�vY���x�䐠��)J;�/8��p �f�[�_��������調0���R��?a�+�Q�����թ/�y`�(�z(�g���մV�(*�`�Xa ��Ea���"��>����$��jW�7�w��:c�S�>ͽiߡ�jF1�X(�h� J������f'|׺�h(�:�I�6vu����,�
~�.G�Szv��� �,�[�;M�~X���TCD�(x�1��Y�cޤ��ŵ'5IP#���Q�,b�(�o�T�[��c|Y�o��� ��2���b���S�>��� o+������NB+ G����=wl_��n���"���-V�D�>k�8F��ę,� ױWQ����iL��~u�+��H���H�F��
�#�j��J��C�w]��8N��/=e�pEg���� d#].'fX�/���m�SV���ǲB8�"��P)��Ch�	��ł���+y�0��w9�<t6\������Y�N�0�����]��IC��t�J8�>6�7�8�V���{���}>:h%���㒔�I�eVzٺx�:]�Od���G	qƜ�ٯ�w�wC!���s����)�>�,T��Q��9D����x��5��4���q��!w���snk.�$.��M��v��d�Y5��};�BX���!86d���Ոw�L	�w��	���a�X������"p)G��j-�LR�P���-4�@A�*���f�f �� rw�(X���z�:��K������#ڗO��U�j���+c����#!�G�ظ략��5q��:�qÂ*�n�N0ž@ �U����5�<��y�{�3�bd���F%���l ���!.ͱ
}u�� ��_�����}��΋�!S������'�词ן~�K�P�j�+vZ���y� ��1LT~��J�hr��ٲ8�T��V4-\8)�W�5�x���8d�:7����П�&U�ǅ�Q.���4O��F��0
�Ę����G�YZH�?R��ضB!�1��b�gG͛�|l���u"�Xgb"X�g6K�*~[�3�CM��>ũ�%�ƞ��J�����d����B��~N.#	����%�/K�N`�7����y���j0��^͋�,������i���~�����
�����w�Í>Yaw��F�D�L�O��:�;��JJb5�-,ޡ
�z�m�$#E[3�bUO�/��igAq׻����)ڝ|	*��O��x_�;-x�����v���_�%�VX5��D@w��Ye�-��_j	�{�uX�3��`k�y�[��?ߗ�`lu(3}&5��	�C�o�+����R��B��������eoVr�Ԝ��;:��{x�
�j3bJ2�����0	���+��0>d(����P�60��D�E'�{�èl8r��v���#���>|�������
�k���P[�����'�G�[޺����|Ck�/�(���,���]n��l�6�0@��?Ԩ��:8�S��:9�r�������U����ڳu�38�}�o���������~�af�Փ4҂7i�Ҳ��|DE�*�*�s8�z�C�Q�x�!}��q��{)>�_I��$�$�hy���Na��<M������2|~r��AP�\�i.AU;� �aK}�ز�S^T\z�.xr��:����S*���x�|ԏ��D�V�1%���˥��,:�W�:��z�Ti��x���`qR��fEY�/����J}7�	�@��M�xdf����`I��#�j��E_d�#S �<�C���"3��L��V��1�>b5�wFZ��U*bVl.sG��qb�b��`��10�!r,�aG�v�<�:4se�w����'6,�� i&[G�mX@%�����|G�uRx���U����q.V&�*���c�j#�ܒ�Suk�"4���ȟ�T�n'�M�? 9F<ꖸW�{B4O���a M�E+8��	w<N�sy	��w��Ɛ�v��EN��D�w���h����ד[;�b,2�B��{�}��k;�v�W��~6.sWkY':/�G�
���͑�9L�K2�u�ft9�'��rd����{m~�o�Uh�� ��%t��8Hc�o^n�1���[W@�ֺ���t�	�k�UzP�A�,>�����/���P-lS�����ȩ\�Ɣ�U����dJ3.pi�U����������*�cȞ��Wy�n �*Pd�p^d��J�,��c���L�%T o=1V�O�$(�tGe@��R��]����v�|,�t(�	X�SC�x{ �"Sd����{q�I����>��L�T���q>�ǁGʯ�©3����M�P��~b��č�Ө�&Z,�(�u���V�Va����������/�I�Uz��4Y�-�zf����>�X����#"��T����K~h}�>(���$�k!�'�����m|��:x=�>W��Ҿ�q	�|0����	��I�MO����[��c�t�4��s|��S�����O�.沭���j+.��un�D�`���4T�,��]C ��kl�7ߒ��M#u�.�i�oZ�py ����#�5�}�(�d�X�T�"�j��r,��7Sm^GeELgCG�mܥ	�h/N��Z7���e�Q	K[W��Z�~쭸�V��T�,\�#��j�H?�ή�7�FII���������.+^?EA歷�ϋ����O�m�s����c��iG����x[b\��?��Lߑ���1��>"����EE�yd?���>���Y<���D�p�N���3˷ $^O���p!��lt��|{����z!נ����0س�͒ޓ����|�	~���&�=$��%��7�2�P��K$��]�]��@?����t���]�G�x�%�����з�����`;��� �:C��K�k�O��}�d���r�
G��(jq�����kK��/H�Y+��[�F�@�A`/U0�1�~a�k��S~n�D�aع���e��v<�Q�����(��qu�2�F]"͟0U��I�mǔ�C�Q�*�ԥ2�KӅ�-ro��a�Q�u��5�6s�*ܥ�8	F��I�9&��W���g��x����t��Mpn'�I:ϣ.�.����~,x�@d��зz-� �^��sg�"H'�?��v+WP@۲Q���Ϯ�ۄ�:���'��2P�QT��@�������r����� 9��g�����k�4�4-�o���ǂo�#|��L��lZ���о��l-:3�gɏ&���o�Û�ˤ;q:�K?�Y���2ͭ�l|K����iY�Vvpτ�X*�z(�\f�m�sz�uF�'[&�3. �}&��H����y^�q\p�ꞎ3�� '�K��*Ѵl�́�}|�͏ك
O�\����O]�4>L�t'2�y����V�Ӹ�_<Y����������6o��ˮ��
�pp��\q���*�'^
t�o����u�i:=��y�7H\ŅW�[Z!s$���U<D�+)���U�}r�obhH��.�gэʸč�x�q��$7�t��
7tݽ��}�������L%�CrW�o�p^�?N���/��lM��m5�<y��J^� %J�]y� � h������a��pT'�j�
;�p����ED$H�3��%��g�攩{L�/�v�Q�!@.�'���-�T3�K���z��Ԝ�;=�)�5zc%��j)'Ǆ "��pc��@�B��R���Kq�nbn@��"�n<���pŖ�9�5@X��EC���$J���gj�U�I<YC��.4�k��
�c�yp�iJg�mL�}�g	��__+��㕰7��C���i���6��??:�xAD[y���9��I���̓�;�]��d���:dX��"��٫��,ʨ
�)L6��Nܩ4ZT!cN/��X�4��̸�dYu�DG�y��?A��k89�T �i����$�o�6J������b�,#��^q|�s���!���6������Jj)�-i�NK1�w)ꟌW%D��ݜ� ��'5�ź������M�"x�H;9�Ρ=ΌsGjGf������_��;������8.���X&8m��H	��SwUq�o��/�71vު��4J�Jr�E{H6���;�����$�+�pb�7R�� i;i ��'T����ީIJ���s���l7����󦜜 ���I�@kS�N�jχ±6み#i�G��r<�]�G��-l�*/�Av�+�q��c*_t�,u�-Ro'O������5�s$S�A~-|�������O�
Z&6���RxF)y!�VU�;Gñz"d������g��`���Q
�#���csh��%�a�y3�z_�Sn�� �~^0@�'��&�|H���c�4�o���~��y[��A0o�`���=RD}�b4��KKi�	��+k�"����%�d��ώ�45������ڝ�[�Eh�q}���a)=c��hh��Y�km��Q�8~@IY�R1� 	��,�,�]��� 8)-T�BJ�c��z�mE5��4vt���r��dr9<���2M�~O�g����h-���b���15ѽ�mm�D�{TA����B�N~P_6���@JXN�حW��ZÐ���<Y�,/�twOA���JyV\ьتO[b�E`j�ROWqQV���X��!���V�V�����?AH��v�z��z2�i�O�����:�[�nĥ�/?)ƾ��Df�a�1�[����	;��b�2�ñ'L�)G�l�Ç��#_<ܣ G����&<l��#�k(J��E��%b�5���d�S".�/�����Һ���z��.X�� /�zJ���"�G-2Ղĥ��w����n=�5����j��K�a�c?����A˫�=��~����U����JYe�+�2�Z�O|�KM��3�b!l;��J��X;�����kDp-ў�a�����B. ���T��0�9i�4a9_=��+d�~�;l	��a��e���{P�!Y�+:|�N� ��D/���ݘ��̋���_��l��i����3b�b�KQԠ���P�7�9�Ian<*�� ~�z���I�����D<aQ���6P�]p|�o℠V���aA���K����`�;��ϖa�F���1�9&��y8��4��̭"}l����ޮ�E��ܙ;���
������l��l]~4��[�@ǐuy$3��-�7�_��5m��wXA�U8� ������0kN���p+�U�|T��-mޮYt��@�uINH�1S��0Z�Qq���Lhd�Ɣ�2��M���~�������D�K��"=�n?��]� y}����r�UǒY�{��vI�l��lC�;����3��<Ub��Y�4=�iC���)p�����qq����R�1#BW�4_17�L�
5���:C�h0 |������<��0@��'X�T����� B���-eI<�\��?}|����u���i�Ab>ϔ�2���h��K���ve��(�UbD��ӹ={-ʳY7"��wW�-%�,uC-��:�S�<�s��f���s�^i)�Gz��W��B���E������lt�: ���7����z���7S4���*nN�롾�b6$�l�N1��cŻ�6��o׀�ȢS��ք+g���}��^��"��6e�K�[tBc�_e�ۂD�~Oz��D%q���3!�v:�o7�Z�7k
�8��W#L��k2�jU��K��[��������e��PWT8����]�?/��l��)Y��}��'�o8	�����W5T��Y/�ROg�b�06����l��1q�[t޻�\����Rv�멯E�PAT��+��	�w^��Y5B p�0���r����	��a��e��f,�s��Q��3����OUT)�C�n�k�� \�z���9s�t.!���[��rY����Z��|�$ԦjE,n�g�ረ�L�8�=[���4?��Q�%�%"�擄�RΏ�[}�3�/�,��t_��1���9+G���{�{� W��9z�0�9���Na����(�B��#o�9=d��p���Z�������5������d<��7	� +���K��l+�d��Z�x�yPǐ�/{Fm�VJG��������a�'jl/'��Y��{�f�vO����'m@����d���!�=u)*�`3;�f�_�f�r�����ϸ�}
�:M�H-_x��e�|�������D�<�	~�U^e\6�S���#�2tv�b���..����'�������VM�!A����m4�eoi�����ԭ��!�d/��`�R�j)�����z�����)@N��T�m:�%��z+�Gp��1��##�4Į���i�ZZWB2�C���V����`Kv9*�Xv���x�q87��O`��_�MH�Ц���&%�kgZգ^���w�\i	~�upv75���j
 I�d�`ƭs�Ѽª{Û�|�����7�������\�;rl*QQqr[�<�Y�"e��tE�H��,>Y"�.r�T��9밗�+�dXI��?��j3�!{�������<X�n���疊���5A}de�¹���C�p�2p_�ƃBN@7��K���c�.T�`0��T dՠ`㨝�ȳ8ږ4�D���	��1��B,5+磱-��hY���>��Y��}�����)�A{.�8nÄknZ���)5 D���JCk_شl��tI�3�s���X����{�b�@�(ocJ`q�
��I�2VG���������J�Q�U����|�����<T�B�`"*�e��cw�z�`A��{pm�Kj����sY��?#h���;Y������J&�!eQ�	 Y��B����AadBtt3Ix������ٔ�-$i�����1�2�|�����N~�Q;l���suDԉ�<���"�M���W,��ЇD���\�>�0�p�� ���nǌ��L��$	,���θ,	�T��XK"��b�x#F�q��
P����ӊK��G���U����x�TsE��c#Ŭd�0���,��G/�$otnWo��x�F +5���p�6����y%v�r����B�� �oc|BVo��ǭ�ϕiKo`�W�Wƴ��sN�ԏ�u�A��h�9�aW�P�s^ZQQ5ZŘwC������L[���c}�����3�-����|��e@�X���|�7�T	pӹ$t�±Z��_�tu��
��ᱽ��J�����9w��������KǤ��s�U�N��Ƚ�U�}H�93��/ā_q��!�%�f�B� y�KXk"���$�X�oj�Q� �4982���,_9g���j ,���s�j�@�c���J����W��	%�I:��6�|:��?�Y��*���Cs���kMt�>
;��W��R��Q�+!���W�}��6Q�Q=hu����n		ZZ��c�:!��&��'C�4E�\hg� �����0I8,kh�imj�	�t����������ɵ�+O&S�kO�қ#SN�c~2&:�Qb��OT	������5e!��~�X��:[�T�P-���g�4����Pr�b����(��ڤϲ����+>�n��k�Pc>7�Lj[n�7�T�n7�U��?����Y �
\u�N�d��sӍ�#ײpO���t�����]�5;��O.�<n��C�pnC)��֥���T�[�"P@aox8�Mߓ���}�����=vֱJ��؄3|afT�^�������#j�t�>����P��4Մ�z(3�S��a9�.~����Bͥ����(������e�p0�5�V� 4[B��v��I�Y	�['
ͤT��$3{��~몙�ц�cH��#%���0Ǆ�a/���h+o�����N���?�
���9	�Fߘ7q�g�D��_�zή�u)�����Q0b-14�_�����=iQE9��Di�<WZk��/!�х�
��a-��锈n�:�īz$9��z�F��)#�����o�!�M~����)kA�,IU�k2��L-b	K�*X�*T��4�;y�X�k�7}*B����뤝�y
� �c�D˞�h��s�'�E.VW�6�w����9�,�`qG�,���WS���8�en�w�ہ��l�>���sъ�����1}r3yN� 0fE�w��6���S"O_�{����+��G���rj��@qĖ��IP��ujR~��\����lZ0�I�:��V7� ��jTdZ�G��Z=���"��IY1���t�|Q�H~5&>{�?M�c�����-��>�QBD{VI���c�47��r��� {��]'#ߎ9���HG�{~�y�<ղ�t;���M���?LW�&�~qƮ��6`1�k;���A��{��՛!�w;N��:��ғ�>���b)��er�ɞ���
���H_��w�)Z�C��e�G����
��8��#-N�v�zO�/�ѽ���߸�Q��'�>X�0Ap��-5c�R=d��t4��h�t�� �˙�-��Y�Gz��aM���CY�{��I�.�j��+�TRf�+��o�x�~6���O,�'�kjO���qU &HM��R��S\ZV�h�/�.�d�&sG�w��|�W�|ICj{��p�Q�3\V����{L�Bi���;��'>-�%�yzx����Xv���R@F�\�ǚ"|�!�{;�Tm����oM�͌���E��&�l�I-yj#��$� ��&����lX��6l��F��a>�v6�O�0�|�IMX?�6�o�x�Nя~�z��_a��5�Y3�wh�yJ�3��2$��u��+S����I3�i�<ڔ��3��UC�*��R��T�$���ƾ/-��[ndo���1 ���i⓭�[ ���j�Qe��e0���QZ�P3BT�"f�c�0rX�F�Qy�݋Cd��8jY��-K/��W�M5l���vO���ձ�j3%io�N�P����ނq�#����פ���$�jY����Lk��S���t���t5�)~9"0D�����ڸ�ny2��Q6Gjd>p�7~��
Y�RlF.�yɣE$Irn��rrge����d�:E��I���E�ȍ[�惰��1�p�K�a� ��_c�`X┅<�33^�+�ygb��zz�¹e�( �'�g���&��S��1[�1)�7y*�ˢLM�)�'^�4`�:�D�[�Hb˲Ch���S�19졯d
���]��Q�-��ϻ��Y���� ������'G'h����\��aW���C\�)	�2�ȋі��4Y��F�+�kE�/-%Fc	��L	�~�쭄΢`ӆ��4MD�yva�x�>�bdq��I�R?:��qN��i�oI�5FS���ڒ4�^�K�D�A����/�4]|�6����,����%Y��z�KU�v����#��釜ؾ7B�{���~n黅����x4�Q�\~���+꧎AI)J,:���l�P���5���'Qv�*��Ř���ο>��v��k��c6`ں��i��}�_eJKFTS���ύ؃�q+��R�գ���s���z6
p�6�-���W�$���:�T��4�v�E�z`A�n������os@�ZW�u�.�ԍ1���M{GtX�V��D)�4�=1icu4�2Z<hlY��[�	�������f�rЋ�2L�kL~��	wc���jh��n��,PK҇l�,QX�;��������&����S[?�i<�2�����20R�z{`�/f�FjmPG,���e�������r��>|� @9m>��K,`WЭr:����~ޫ���:���#6� �N1W�`<q{u7��"J��9E��^x2-#6L�J�]��IL+��P�WL/��[���2+�|'a|�j�M!�,9 �D��~2�����~��H��'�."��+��fTA�����Y��k'v�OQ�s_�����Gy����ؘj���eOtZ;HBG7�� ���B�ѕ'���;�ҡ��Y���>'�f�m\\N�ͼv������	��*ρǼ���:����߅E`�sx��7�B�j�2�[�ԼVj��8}K��H�e��e
�G�?�@Z�����xX!�ć5�����w��7bRZN�ڍ�C#��,p	$�Z��Ԅ~Q��:G��y,�5^d���#���d4CMBh�nI��,	�k�I�_�bSb2'Y%O��X���"�X�tЇ��A��f�w�p6�°���k�!)�L=�Y�
Gm��Лr!*A�ՇX���� ��rJ�63�`�����H�1��|�].��[|���vY����>q�p��Q���˪`{��B�sEж��k�k��,H���3@t^O���������]&,|������!+��a.\�Y 9���k_���jS�
"�Ɛ]���R/=�j���/8뭘bG�l2
Ho�K�|¼GT1����X������}gn0!y
��
��� 	.Gn�J4!�?�WG�r�nox�$pT��Y�]�C�.C�լ�,)В���aҩ��C]�~��Z�����?ކc�Qn��|Ϟ]�O������	�	���=��(���
�FQ,�e��eEC��5m!]X�+�`[k޲Г�����s:MktA��ru��#�ɧ�uU�t�g�{�a���ʲw�-�:��4����'��Y��
'�����X�H�0��v��9���b�Q�$L�	d���\8� ��%����6J��z��8f=�|���g���yvD��ټ]�]C��������K�Wl\
���ɔ��/.;(J��;	�̾�I�1�������4�-��G��ƕ5��m<��"Z�D�Hع�sH�d� ,w˺�c����[��D��<�<&���F@^b�˩�H�FF�?�E�� @W��CN.�����ʫ{�0)5�k���v��(�_���@��A�y�m���֔Sw���p��2� ;x�`����B�;�\$����DKJ��vc [K��(S�(W���N({+�e*x�����0��g�ኜ_�i��_&�h��N��|B\�7�'|a�6�K_��(�@9�O���4����Z�~aI�w�H|߀ф�/��]�u�Ļ�iG�����&�?gR-'2�F�Zރ�������s���X����hSkEum����0��ls�e�	�Y�g��/VK���㑖����B僧�n<Qwo�`1� E�/O#D�e�4���9!���D�)�ґje�~�{����q������ ϴ�)�Ł�':��γ9"8�e��
;a����3�Rʷ����L�/���K��خ(W��	�57�?�p�A� +_�`Y�W��<�^+3QDQ6l�~Y�gѿ|ʂIO'�0��O.��O
�~J�,�9���Y5����ců1N-�:�{E�_����L	�!��A�>��Z���p�ҽ������]�8F��$^V�
m��a[.�&Sm��� �q� {H��W�kٲł��Có �!gɢ��� �J�?��/������6��-�d��R>�Q\+"��n�������@��gy�<ݡ=Fy��P�� �� �ћ\���N���Jp��8�w��l!�~���Elm���\��WJ �S��p�aW�`��W�
 (`��,G��,R��ʿ1�[�q)/߳�-���v�]�Ź!=[µ�$�S��z�#��MɿI-)m� 7��?Î��^��P��'Hs˓�����@�6�4,��/���,[W6H���yMg0d��6Q޶�]�K	^�|(��wT���%������>J���F�fώ�3;?��b��O��\0<E���-�^2��U�^���,'���g�,�oR�/��MIԢ1iS��I��@qEL���[�K�w���K5w���{�U`���\��n��A�c�{LE�o����\$>M���P���r�EM~�������٣�@�;1{	Aͤ���=\��4�Ǟ��K�����y�����YF���G�6*Ff�K{� 7�GF�������㎢bc ��6?����T��	�>P6
�"_�K��JZ�(ܘ�`�W�d��߾4q��Ԑ&�P3�3%K��Ԛ{�Os�Y)���>�d��e%�花��?|�G����+����Й{/����{雙S�|᜻� $��zոQp,�u��%[H�z :�0��!�"�"h���u���r�5��}�o]d�LlE��y,;&�k� ���'l���0�X��`[<1�%'�:h��{	�-ͯ%'����Q�H:f������4��-Z��S!R�{�}E��X$��2K��<�d���_��x�j����|yI��V���|���mg�lOd��� t�����^���#=ٚв,-׽H?@d�8�i��h%�ci��H�W�ޓU5y~)E�?�{��Bcb�q���m��?���4����G����h
���ԣ��ϙ�q�����+�N7]�?�'�-?KЁ�!��ʇ��SN�@��oA���;��c���� 4���fz`����5(C5#\�� ����߽.u�>
D|y�-.���}b�C�t�
�C�������:x�(ثv���_�ǁ c�9H���`�R��>O�9�P���B�g�
���2O��S�P���:H,}1�BXN��1��,��l�9��,�4x��*�S�[F�GZ�[];U:~��,�6�,.���1�4���(T�A���v����#��u_�Y?�u�����or�D4�`����lRf��S�Z�r��{yofߑ��$ 
n���u�B^�t�� ��I�C���2�s���j�m^�����U�˶����4��\֊]���q��X9���)scAG>��.�6�}��~�T�E�k��|=˧�_=`�p@��<�sΊ�Ab՟E��._���ʐ&��zȼ��F�hn�����+c��x�����U7����˜+)6r$ixA6Ehp~ׂZB��w�]�ng�3��
���}O�?#׽R��
�PF�=1A;Ĉa��3o4k�Gx�m�B��(I�v���<�y�ɝ�*Ta�T`I�U���N�`V0�4P�r�CsBFɁ���)���VθcW��I<�����A�P^�.I2��z�j���B�'�,��N�\�e�^�o�vY����	�\U�|��J�zĞ��2��Sn6�5�gX@dp��h��c���0�!�?Y
��pP*�ä�8�7��"Lp��N"e�5�='~߲?������OA�7�Wv|�wS���9b֬w&$|�ǆ�� S����kj��	�^��u'�Ov�b�si���!rAy�0e���L!�EYp�R��v!��'G�V�p�3m<Q�M��!iħ�|o�`�㨯�ڱ?����=�p�D�ͯX:��p��9�Ǝ���_�1�:ϙ�� Oכ�G*�>���޻�eEp1�CC+^q���!���PI�T�I|�����L-�d�����������?�U*;��=��f�}~̯�4�׭�Mt!N��w��}[u�;tǻ��g��@x���v�yp���@�0��Ν�i���T�Iq�;A�R����&J`:v#���,SԺj��a-l��E�=� ������c�2GB���,M��Yʖ mx�&��M�tх�)"��U��YT�(��-j�WX�R��M�����Fc�
�gԕ+(��_�	m�\�L�34����Nɪ'L�E�9u�uAa���|>� LɪR7�5�v���<�����k���
��Yϒ՞���
��� hfC��EA&=.%�d5�
p	w��h%<'��j�2=���d�b��v���ڈ����Z�_q5n����)]Hg�l1�B����B m��!'���p@��U���+���K)�%-�>I�뾈���2�?��o���O��i@��V�i4�K5��V�l��!Uhǟ��%&=e�t�A�&J.b�_��`��@�na��掩
X^����l�D�ZC]h�<wt�{�LK�~���N~J�Eũ��EytK����x����:�I��D�d�?/s.���c8�҄��f@8�	��|��Z�c�2�້��M�=�`	`/&��y6i76HUM��Mx���d�L�me�������u���QW�u�ȮL��L<��V�ڇ=�(��CO�4<��T'��b�=���$�����m�!$����s����r 8��=���w%D��BJ�f��`/Ay����|YאQ>����T�ˁ}��)��UGu�`7};�4��2�>T�����T�|�FCވE�L����1]ʟn�^&�礜ٜ��i��Ԫ�����#�V�RԳ�ZZ�!~��W�.xs�2UE_Ms�wʈǴ�����f�ip��7�E�!/u�!�ԫ�_R�qHO|���~���h�$�@�e�X��N� �CpB����@���q־r�O���	���ԍ����xj�7�5�v�ކ�-���}gO:r��!�!��[��d��>7�z�-��Z����5���-�g2x;�`�P�Ə�Ng���b"�^��E���#����V�?kP��.��x���I���L�nx�o.�|��ʩR�z�oi$3���c����5B髎3|�5�N��֡y�ޛ�t�ΐ�x���8=|��q�TS'T�9N�v���U�N�''�'�-Ǜ?X�w� �[����3<�t r��o/��6�f�m�ڹzvv]�˱C�
U�?t�fE��#~Se<	����]�����Hχ�h���a"2Dߨ�(Ż��H*�dU]������$�XJ��P��0��
2H�|KL+
%h4=R��o�h��i!��qV��8ˀ�����A����=5�p@"�[�6��Ʈ`1x�5����b�WL-�67X��M�V���2;�S�x����pꦒ���?_X�x ��'O���A��)��B�e5�#\.��:��M	�i�D�bgIj��	yf8�o��vV��'6��&�&�B���JA��7�
�^���������$�?�PD;Z�;Hn)H��.#����e����+^�`2��(�)�gX�AwZ��	EK��˲�-�l{p��Q�oqD��)�L^�#��b��͎pYsc���㆟gj����մ�"׮�{�q���+hTc�DO�ҝ9��	�bh�+�J��C*��ꨊə!��`��;�~�s���y�~��Y�E��g��\� ���<�f��8m�K����vW�Sa-TM1���fWވ�V؋�kŉ�[iS&i�ۇ9[Vf&}��	fQ;�h[��{�+{"��}�j"!\$c��*��6iqj�:0ږQ!Fº]��"��_ڙ&�5���YK>��=��?I��O���s��A\�3�J����y��V��׉��&�T�ܨgn� '��_��oW����0�6$�����a B<�PI��(4.���U&#�1Y��R����`�Z��m6pw�+2���.G
Be���'�ĒXh��s@�t]����&Br��[9)��2}�F ���oDe� � q��t14��-���)��3�WJ��l#��*桰�m`$�v�k���!-{\�uY�T��9���M}��,����B�Y~Z�(��ja$P,%�NV���w�Ć�p�P���k�i��>�;b��]^������[)�'Ox�QR�Ɇ��s�	�;���Oy-!a\STx%�:� �S=�=ނ5�eu�F�b�4fF�����)=(|��:A�
tq�#v�`Q�ӫYEN[%!�����>�8��n�L�����s���Y�,�qܘ�/,�\o�e��R�U@g�<jj��=��������1`O��PY`ɜL�Ҳ��\A�Z�
+p%�&@�;f�W��l�R���c�L5���'�/;o���1�#
z`���b�e����z�.j^��׾�BJ)�_z޾A���3.���1yـ�����t= ���ʽ���@�Z���N�<!f<��r�M �άl'�8x�p�5���W���3h\71c���v�2W�U��N��u�
C�ћ�B)�2�Oz��^��F�FV�����מ֧sA`���������
6�`������~��W6�Ŗ?$���o��v�1�<Q ���-�hO����D�����h�1���
��~�����~\��wH37�Zh�3�@Գ���&�G��g�Ԓ �H}�$P��	8��?��'���:`�>��$���|��w[�`��F���ј�t�"�t8�� ,LL�}ح�"Ae��,@���K<:.�"�D�7E\��i�����Vi�|V�W=�#��mbL6/��nn��ݚƊy��T熬C�� }ǝ��H*����(�dF2�w�x�5ּm���R�|#�G(�o��|�	rbnA��6���v�L���9���(�biկy�:�X��u\�crc�[��� \'Y���
d� �F�k�ݲq#���'e�&���>�򫼂�?���X?�oQ��0M�p�h#j_�.\6��Âb�����ǽ�Lh��jk�}՞m�*���^�C=�+|ƛ�Nz�T��������G�I�$��R�fhI<`$���&� J����T�I��W|\5]_���]B����������`�=��b���t����Ԉ#73��9��[�A�(�������g��1����F��������X����Q��ҁ�NU4S����2�����C�9�*$�Ϸ[�Vꊑ�]�j���2M#Ph�-M���e�
&#�E��QH�RB���6=���t�� L��bk23yF��	(�BK*[C����h�{]G3�S����P�4�����8!^�28׵<"Ww7{��.����F@���6W�k��Y<��D�;��G=$@����?�cH@��C�P��;º��Ȕ�@WgoͯŘ�ƥ�uj�jxf%���`EvՙX��'U��  OLqmd$V[ᖄ�&{B���-BD� BI,B�^���pe�P�� ���v��@�=a�]��F��uz>�A\��q�O}�d�1c�����������9f�ƿ���2�)n����kTPR;a����7�ķ�OV��~i���(�_uY�EY�eaD�*k��m����b�'v����/0���G�.
���>�����[����5�D�>*ַ�>+Sh
�q�J?�ݢ,v�j6w���cS2�������ε�09��$7:DP�$[�D��,&{�1V�0���зS� �D���[$��N�gs�I���!	�S����(��S�#���*C%*1�������'>����D�X,��}�6�7��B`��\�T�������'���˓�$�-�{���*םO[���pG���U�H�TN�(߰NbEH�u��A_��T]��!a��+�:�Y��Ɩ͖|Ƹ;k�,	�O3u�[|����y�X�YLq�ˏ*+����
��G%�(�,m䝎't�h�;��CZ�Ԅ�W^�z��w䱾�0SX��������_�_BA�l2�.��&,Fߎ�i���$_�0�L}7{���`�H�j���|�	��(��W�矉�;�)�}����Q��D��\��A�]��n�w��4JH�[�r�S�/�:�u����tW&ao^�����D�_;7������#/�	��2���2hίN�@D��X�N��V�1�G%��7?8%������(�2�b��b�k~�������<�ڗ�MC �o9�ؗ���/x�������=ь���μ�!�$�n�T�u�=�uW<�i�P��u_v3��<��� U��٧�o3���N��� �f�1��뻼]%!�Ĉ�N��������(��%F�+a@�~�A*c�?����VQ(D�1[>���W�.�C,̳�H��A�ۍ7�x�� ��>Sx�W�W?���d�L�jW���(3|ïI� }`�������c����.p&F��e%�������Š�����\���T��z�1՞]�8�e^�|�}���r�X��@�c�CY�֪e?�Qm*�q���˸ �h�G�M�,��#DeB܎�/�y�.���*}`&oVIp���I�<�moBM�Df�q�[��&�	�3Ua��Y/��U����ᶶ�j" ��Ɍ���#�P�43�x�έ�*&og$(���@�v(�)-�t�I/2�٨�Z�w�����6�10!�eab���7Ҁڠ�������K�P�n9!L��(��z���Y{3�J7�=��(�_z��s��E�Cr�{������mo	G_�$ �u6zG03+�K'�0�-�6x|�$���S(�=���=�Ʒ��r>	�� ho)"�n6Nc%]��j��'π�Xr�*�Z}�nK&)gj^���]��/��� �r��ƹ/��hu�j��D}I�`��zg#w?U;C˯ZDH/X���AQcu�I�r!F�(�X"�β�ގ$|��g���$�Ib�.H�{����CJ�B��0T��6v��ThƲ[�1k
b7����Cl�S��q��;�=�83Z��b����?�:O�y�)d�����㊯� wp���^��?<\���t�<����	���%S�ηB�a�[��x�d��+>&��t�ƙ|%�{��ۙ5ri~�*:�}ԭ��2���T��{��	[1��L��%����
�Y4{:���Z�^�ܤ m=lP�ض�N1�*3����#+�t�G?�}�'�>�a@�d���J�\3K���U��M,F{v�	5m��e�a���ړ۵��e�R��I�+��*������R�k����t%�qQ�p���Y;���$����]���걑g�x�Y�V(:W2CQ�.�V�)x�cH7Z�s��[X)ɫ��"c���!�lx�&� ZG6�U�>�;q�����[(���$��z�H@#u��A�1�s�S���96��ʛ�����eP<Y�p\�V��Z���s ђf����ᨿ�?P���k��f�D�To��_R�VIJ�k ��������FA2	q�@�ƥ�Vb�h�^�.�� t��I��b���t���L;�I��A�"#�-J/�z�X��a{�B؜��C�Y��H��
~�-�.�*�(��Z� �S�E��K��et�&�!ζ�n�
8���M��u`���]��T�A����T��*L`��3S�����)�X\��bЂ�b��@0:l*K�O��V�R�ڥ�[a������jl�O�3���IA���eՕ!iUU������L���$��ݱi�O}!ڽE[�̲�����C!������aNj���ٗ���ps{��No�%<c�!��kD�� Φ*Ex���"S)��UBB���{ЬVJ�偟κuH����J�5����E�%���S'S����-����s�0k)����專.8 ��QW�I!���3XR{��9�`)�Th��)��.ǹi'��<�5P`?��)f��a_�����¯-��8n?� ����z䥕�����(y��(��!�Ԋ��o���� �*PGk�E0�D�b��6��2������o�[[�=2kז�<e����>ц��+W�����8�>َ��F����`0��uFM��m���jj&Pի�x��T\���3Ȑ�� I���s���.|��>��G,�`�/t��&��l:p8�K�CX��>oy�m�]N֥��'�:���S!#l���X����L}1/;l���j��^uZ��WE�M|��Q8��_0� �
/n��`�% �.1����q�n\�F6�M��:9Ӵ�a�Sw(��*@��휀C��ڮr�; k�}�����S6��J(Y�U�WPC�f���M�NA�<r��������}� *\
�+�4��V&k�d0�&r�'t;�m}����9�v�h��uvoe?=�6�T�����8���� ��˓i����dWg�j0��+���?��X����T�qX�(�0!�{��ۜ[G�<���?�
��9LF)�(\��c��Wb-�C �(N9_�'S��|�[2�(=�����lN1Ҏ�����`ʬ7�e���nEPĞJ#ϒq�X]�OA��p��y\��ʏF/�5 l�.�ԁ�bE�MG�A��E��=��t<�\�lXG�]��I���]���Eu�w��Qd{ ;xı	�`�H��#y�?/1~쩔���Od!�H�p���i���߬���ڬ��89p�_R΄���q��`Ǡ{X"�^�jR�H�
�S���Z~������ �$ћ�<���;/ğ�P ����������n��5�7���:dy�J�X�97�1�J*M�8
%AY�S�B�������[A�1�U,8R�@Q�j?g%���M��;����Y�Dޝiy}���`ѓj�ĲXї;n�$_�Y;$�Ç�DϢz�{|�(���[��0������kB��"�m�c�8`�m
��}"7�"���yz��#� ��!�d���� �rD���z�5Һ�F���u�<�t48ݲ^g���\���-9rz=(�>���s�*%y����&�+[�&�QO��@�����WM��q�9�ع�뺬�ѽݕ'��0|�.�¿G�}=������#��sp�G��/�%�;��(^�`����HDP&�m�U��zz��gP�Ju7�|���H��|4�{W�#46�����PT!�b�()m�͠fm�
g2�3xx!r�^�d�X9��	MD2���O�i@y�T7�;=�џm�����py�����0x)�y�}c8�͙�4��
ǆ$��'�����f����._J�r�\��Q7�FLڴ�o�Q�֩y�ڼ�~$�(㹞��w@�=�d���X�N����e�2�O��{5��D ʤs��;v��8hU�QQP���x�t�*3�Zs_����Ě�����FI��i�g��-�j�niTKt�;R��G6�3^�$���$�R
Z�C9����e�	�p��yp��c��^*�]΂Z���h>@c��|���b�cj7���+��]�i�n�~4�$vRd��̟��_}2P3�S3-jv�	�ڰ�>Z����֌O&Q!���9-�=�Jˈ9>b>(^�;#�KP��;sR�ʦp(��н��ѳTˀm%��Wg^����nm���:O��X����x+��Í�08�e�����W����lV�i�4(��_o���a�g��0Ϳal�y.����2��'� ��'?q���ߝ��y��� `���sE�����f�|�?��Ҝ�e����#!q?�g�֘��f��I���F�����Z��\l�P]�����a�1�6J�V�j��;����fH�I_�S����3S����z���ad�k�G,Lb7O@?N��z�r"X��q��.WX��¾��m�i�H���K��O�uzR�w6m6K��b�UOo��q�V�WqNH6��Fu<�j	U� Ў�$�W?j� ���^
��(_��2�
	�<����P���-@��G��!�	
*��p7Om�zKy�w�0G��|�&N�<ȿ�ʽ��������Ȣ�<0 ���������[<-��K��f�v�Ӊ�kd�W� � F�ph��K@lO3�Ք�	�f�:IQ���!��u8:��#��P�rN��,@�OH�ǉ;vi��e)l��)kh/�B�����,l!).��r:`��D��C�6�.�v�؛�NO7���i(-P�+�U��]J��9��>�����@~TTI� �����5~p�R��ڶ7�o}�*U:�d����6O���K�en�\mլg�(�-� ��äߥ�f��\��F2�A�2���Y.I��ғ�L�ǂ���_.W�W�i��e���թ�u%/�_�*{,����ZT�Z��޴���m\�R���dw�Iqq�X���F�@�Tl�<y��� ;rhAđ��� \�S(�O�(������"���u�~؎M(��ke���]�V���q���.�������@q�l	��ڃO�f������nbk��A����ӱ�xy�=��7��ײu���C��K������hy�,
�|+�~�g���J�٣�.)ث
:��G��k/X�H{�=��%=�uQ�(:�g� t���ъ����V��C��)�|õ���cML��IS
F��x��-V�\�ܕ7+H
�� z���{3��	��ggJ�MQ��P�(����4��@q�۶�-���4,�u�*g�u�=t�_��oIH���.J�+�TW��fg��}X¹���NlW�f��(94��)[��3E�ZZR{��T%�9�#�K^ �s�W9-�b�63D?��#���fu.����)QIG�3� a�2����yd��i�e�6?q�?�3��]D�ݤ���y���3�8u�w�yg'}�2�NoHrֽ���0�7�!�8���2��1v��Y���c˯�f.� ��.9��2
���"��٢)�g��	��(�иM��!���x��>a�kZY}�gH\3/8�˺�1�&�G_�g����7D�5��W؄r���t�R��3Q�Q��E��������Z��t����/B~��91�j��zcC�A��]�cq� �s��I��r��c��;��Y���8uDy.���f�����9� A�qz�e3�^��n:B̙��.� �oLht���r�W� �% �X>�}5���5��n0�G�߭��b��"|'?��*�ɢ�J#=.�㭯#\�j��&h`���V:r�j㫦�;r6�f�zVdqLa��%�BN�l�趝����d&ݴ��1�>��L�ƪ	}~TF v����o/��͓'*{g-JW-��J��E�d��OV�J�r��ܐ-�4�� �$�yי�{}�[J)��k)	����-k�k�I������U|��Ӛ���C�ɹK�+�)�W�Y�;���S��к��ȻX5?�ic��y�P����Z@}N+y��>��㶏�B�֖G�� ~��J��#G8�]�Y)^������C���`V��#��@�I��(ڦ���bB�мͣSNt��2�}ᆍk=�kc�J�0�zV�%E���7rF��~V�/�\��&�ק�e"�ݻv�)P��[`N#!���4�?53�	]k<5�:�<`��سg�8��D�|}{K�7
~ޛ؆�,�`�X���wu���q卞p�'L�w
��$�dI��!�Ѻ���CӪe����v�n�i�iB��A-��)4� Z�A ���]ܲ�l��=+�-<|ۖ0/o��KZۇ����
 �p�Y�WܤW�l�`Ә�o
��s��Jk���f����A�^��@��B����b]��m��H��c'8�����^�X2�u8d�_Q�|Z7k  ����xѐ���$�CQJ��jA��U�7��br�ߦ~������'_X��+��X؇��1���l8�g:�о�����x��Ln���j���
 9�m���B�V�*�������}�����S��w7�Vi ��:^آ����xt�F�k�	_k>�7i�I&�Ri�_��:�+>��E����f�ʮtY^�NN}YW�t��q�e�����ۂO�Vfs���6Ȓ����L��[hs�$:�j){m�)�Pi��*����f��b��:P�m|�J�9��+>t�+8� O
�Obлր$¯�L"���5!Q@�Vz��6�`g�Fk>KÕj�O���e�N'�J/�Iu,
=&�?��n�YM\�ӳ��J� �� Hn��.�WBDߑO�E��~���mj)�fl��*���㵵a�\�0=�q<��n����lb��6�Bmx��)0&$��F_5�{?�u�<Z(;��,�9����iT�lP���w������oo"s��ۖ��l��iQt|���;ˠ�x�bacLe�#�w�mqt��4���zgw5�<��R���u����o�I�	VSj�9�:�8��HZ�%�k�� |`���_�~1��}�l�ۧm˰9'�[o=��5{�*�Il/��%����3ϻ8�c��(�kb>��������k�b�>&�l{�@���$1d/���I�W徕�^�A�+l�3+S֔��Vt)�����0���xI}�*�w}��m�^�H��2"P��l�C�K%��k�ղ%�Q/ٸR/s~�	i�mX5.|�J�}��;D�3?��=B,?w#V������i���b�9��["�R���- K�@؊�[��u��{�	W�����i�W��b��1ލ�7{A�����+� !G�t>�It�j����ﵔ���{(ؐ�Ć)�?�pS�LհU����/��=ғ�`l25��~��9������t(r��7D�g~ ��e5§�H"
rqn_����CœU�l`fجt��N���Kg�bVsbma;<f�Em����>k���Fɜ%X#�/�����ѥN!�0�:��*����/|�R�j]���צ-w[K����w�r&�!{~?�9�u�i�L)��g���Ӭ]s�)��O��h��5�E/��-Q�J��d9��-����PSd�ad�#B\ ��Ի��d�L��n%NvuN{�V#!�~mX,Ġ@ݣq\�B�t��p㤶��f�dU�in������l2vL��"�X���}������:�.�g���v�Ql/~�h[�w���F�
�tƢi�h���^�"�q7�x8�P���d��m ��9J����"��ch�ML+��-s#6��b����������>݆4��N����m�H۟���Eo��Na-��֖gn����^�GY�A�:�/��hC�l��;8:2J�q�w=��sh�71U�� �����}���DS�Gz8��]��ޝ���m5���]@ڛ#sVY�Լ�����;����m���gW�x�E<�`�{y�ɭf��r�t��誓�JU?������5Y�UJ�z�I=�b�~*���cD�j�V� �z���2���Eg�g�$=L��@`LG��=)���A�M[��wI��E��7[�~=4��ظm7�^S f�BG�*{
�#mFI���<v��3������
���u�0���u���B1���b� ���gԌ4+�X\� "�GƄ�a}j�,E���7���QN.e�D�R�0r�8,�R^�e��o�3��
}�_�b����,�L�r�sy=W���ﶭ҇,�� i��3�5���e�����n
Å�#��ɫ�i/��>��r	ΟQ&�P}F���p4l>�iD{����
���5����۳
 �}�;?#�5ݭT�-��4�X!�ئ�6��f�>��|_N6�{��We	�}?�ҟD-����;,A�F��qv�gC*����]+�3���Lރ%`i�%+����k��¶х6� h>H"!ѣM� U�)H�r��X�wДaM�e�d�:��] ��{7t&_� R ?���CƉO>\t5QD�@��[��c�5S��ֲ����Q!J�m�#�1GKQ���ی�H߇~������dT��#���c�i_V��ɖuCX`eEU:��C������3$u �ZB2�땨�^X�ob�;���І���L����۽ʨ��fA�Ud�z��9��I�£R���=1�������2��QbaBj9��5���%�^&ۍ��FC�5	_8`���w��l�m0����Y�"76���a�M��<)�p��KT�W�pF�,xjM��'7����Z�өB�?h�S7\.��H�������vj֖s�I(5#�y����Y	腜��V�Mz��4<1���I�(�.s�a"t�p�~7�F���$>�h�0p��Ӕ�]d�Y -�'��{Z�W��j6��g=�4Β��r}� �����(5��+�z�bH�}uP'K�b ������jp�:d��9��J�/+�bz�/%�?0?fp�͟��l����判�v1��]�Z$<�=K/�l� ,N�$C>��X��*T�U�q�	��""wp�����r���<��r��d�w>�i�2\�(A_Y��>�48 0�^.5����2�(����܇�t�Dߜخ���d`!�8���wo�a�F��y�*���pr|�ݬc+�8q��)˞��l�V�P�e2��w��n�k�~��t�v�>��vC�)�:~�g{f�
Q�WA\E�6��N"����e�Iv��5-d�C8���'pC=�v�c�,,�^�O�g~��c�_��kr����G�\����^#a��"�-F r
�N������'Ă�4K��"�W.Z�Ҟ���ɸq����6G�T�����zV�ݸ��:e@���L�/3�}��ȉ̘��ٌ��݂<�#(�TP�b5X����G�;g���Oïc�w���j<�Y���J ЛA�X�UA;�i�JL���C[c�� ��&	$x;xT)��|���Y��!�&Y���ݟ������Q[w	������)HG/7�^R?�n���'��S�s����z��_s���͂#������*] ��F����������e��R�<ƛ<���+'��1�4�9��N�p��\88�7�ȃ�����H��q2=�}���*c��:��s�p�1}P�s�U�A�<v&�����R;D��4�$�,�E�3����	�Ϟ>(��U.� b��I}�$ȁ�9��6ap���N���.~AuU�`��Ǥ�߯���4ݰ��`�� �G�U���wC�Կ⍇GA`��)��B��I�=uQj�ɟ��\S���X_�ļ��<.l��@���E7ؕ��O ��wwsAGH��g)1�����_:Ẅ́�����_?s_�8Y��8IY��y�K����H���d�'�1���G��늵��;��(g�,�d��9���AD5MK��$�Am�Ô��H��%���c����&�ȱ.ꤷp{�DEjεR9�c�'������A6Lžs�h�V9�2:P4�H�\�w[2�!��`�&h�`����X������.��z8�SeE����w��&;r�%��i� �&��O��Dk��/�[cA}�R��myH�j]�<M��Vv�JW_�u�[��#Q���J��ڈ����2h�A����������J�-m�;`���WN����l'�D�J�f6�����i#���_Lt~�<��ϊ���O�#�G��Zk�+�t��mgȎ���J�Q���n�7���U�$�[w�"��ؽ)ٗ\����m!٢�K�����j��'��7���<a;�-h��~���OP<ȇ�F>`-��H<�E����fO�pu����"���ƭz��~_]Vf�
"����� �o��#)2F�4ࠁ�U���a-|���	6���-�;4�lۖ����g*���u^����6�I��R&�:fy��H�@�\���75�sJ�+���Y;P+Kg�A���)5��贽=�ɤ���H��h͛p�N�S�t�߻�����g;R�@
 ]� ��W��^7B�5�AT=I��p8���Yx���e�ԏH��g{$9r��UV%�����L�Sl�� ���pE��7��p%��&�a���^�2o~���^��T*�%7~�ܵ��@�[����*��nA0v���s��)q��*�<f��յȔn� ������$1piF����v�	�Eh��J}{��T��^���Γ�9#CL�qRϪ�ҳ)hQn���Z�|��������p��B<f����J`����e�����؆$𦒦}�XOyW��D.���j���I�N�TKIPt��yڤe�m�_F�^OUBm/�-7	NQ���]6����mRY�.������L��AEH����`"n����9�mk�ꔲ�;��`u�#��}@E��	�����_�e%��J��V��V�D�k)�T��YZ�}0q&��bX�oBVݨ��m���Vf3�cj���sNf�G׽wT�΋��_�q g�o�aL)�B׉BR@��r=�v1<�-}C��d>�����)�jn��!�#F��fs��Az-��a�����_��f��R�j#ő�?t��[G��4A��?9;R���x����)1j%a�&Q��;Y���Z�k�S/|�]c��N==�ݮ$P�k f��G�oi�z��>/ٰ֗�v��@!GR�-Dٮic`	��&=�?��ğ-CE���2~lA�&m�\�"6�*��C����d��c3�S�P:�aMq|�*�(�V���"|k�5����W�YGQ)�Pʼ#{�ªW{���7�E�ZL%��1�a�xPp90y�b�1�7OK��Amw�`�N�؝�	U�	]J|�2V�Xiȋ8�L�$��2\�W��e-�w�-����Wz�hiL���j��j�_^��&)����D��u��t�%��.��\�7s��r���Al�w�24��1vd� ߩ�e�g�1�,�GA�J��1�Z]�8�����0q#��Π�������H�?����$R��飳��F%�	ִ����e1?�&GI��D�u��𰡳m����沟jU��-J�r��;���^,Kf𧽄�b@�)��&�0|������w�7���p�������|{k��T]�|�x�$�ʑ�¶4=b�E�3]Zِ�¢��x^�G�T��*��2�cL+mz�Ih�a�6rp��SPܠ9����R��.���^5�ˌ�W{�B���GE��`���Ⱥ�)�}r<`��ʡ%Te�w�t6Z��Hb�$�%!��I��{ � ~��Zn��>����_y®�����o";�p���d�=i�u$_���{�3������~��+�?-�����$l�r�T�`�����c�w�O:&��_���(�{3��r���x4]F�iX�>�-�\�.�ֽ���k����
���~�o�ePaoQ��a��:SU�7�@{4�ky`_��U˙R]\�"�5|@����'��=F�3.�����T��"�&�R�aLp�Ӈ�^�І�@�-�0�؄<��(R&���u�QX_i�+7�0 {��A�||!=��Կ�?:��f�p~��'�F�%B�r�+�h�ֺފ�g���mޡ�bsk�w�(�w��`�.�E浴J5�&��P���}��[��3��Z!�d��[C�M�}��C��Z���C�?�E�n�$Б<���C�!(}�������n���z\�|p-�zز��(�'�� (Kv��I
r����El�AA;���5��z8�0�c]I�W=9��1ܖ��Y�����ڈ����/K�m�ۓ��؎�� ��hw)�wdf6hi�ʢ�����؜Q�Ľ�6���y[Ӕ�W>����Mq1������_jT��c�����ts�(��Y�ʴ6��ܖ�N �[�6ޢYF�f�b��reӂ���DI�� c�JP ��q�ON˺�,��(�?��XC�8Lx_�fi���O�W�g���}Ő�M�,%%��⊏c�M��w�d�ԟf;�a�����G�'�ӊ䂨���&�b�oR(���rl�GE�`�`NB`d�v	x⭳ǧj�����V�Ƶ��;�~��h鼓�Ǘ'W{)�wb/�zt+�8?�,�q��c�'���\�f�0yg��cI��A���~n{�]�h�U�mr��C�XN�`���+n�����_#��i���9TWj&�K��e����l�O�����`䍯^��0���JQ�p%��M��.|�s��E�?]���>d<A�0�������˓8(���~�$:�@G/ Yȯ���,�fig�
�q4sR�x�(�$x�����W�Jy��� K���<���m��dnѱ������׬�H�� -4�kxb��Ĩ[DW��$�0�3��cO��I��	X����Ոӷ�YN����MO�C�X�z̥���������@�4�WWv�����Ѕ�׻d+I����#W{�Ƶ��A��i�⟙q�JE(I6"T�c'o��Ƶ��c-�@�]�>��>Ѭ�m:����J��r����
�7�6��9�-�-��BRv�M�Y�AꎺY*ᡞ
�Z�0Z�d���R���,4�x?�wIDm�5gˮ��x�w9�,:�)�ЍIx�5�0��.󤚫&�I^2�<�?�}�$�_�����#�S��i#F-C�������%A��R?2a[���9{��n�J��������I�V�9�X�v��ژ�p-p��T�����m�A(֏$]��O��5����K		����޹F,�`i��
$�ar�B��~-�n�65Ol�V��e������ו��O^�:<�nc� �2�'�kۄ�Tز264s��-��z�"�5n)&�<�����8�%N$����q�$���IUu>d�>ؼZw'���pk�u18��BC�����d�F#
���E�
Y-�L�-�,��X�M�b���܆	�C��N����n��U��
Û~q�]������;	+.��5��c�v,,���k���/c��;\����cW�H��0�h.v�:3]]�N!�,;̟Zm \<��E��;��JJ+#x�4�ԨH�1$b��eX7AW��[�f)��w��������D�f�����Ĕ��eL�?׮l�D$�<��m,U��W��훔,���H��	 M/*I�vt*��l;ub@